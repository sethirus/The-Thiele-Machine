(** =========================================================================
    ADMISSIBILITY - Physical Realizability Constraints
    =========================================================================
    
    Defines which Thiele Machine traces correspond to physically realizable
    evolutions. This is where we encode "the laws of physics" as constraints
    on admissible state transitions.
    
    CRITICAL: Admissibility ≠ mathematical consistency. A trace can be
    mathematically valid but physically inadmissible.
    
    ========================================================================= *)

From Coq Require Import List ZArith Lia Bool.
Import ListNotations.
Local Open Scope Z_scope.

Require Import ThieleMachine.BlindSighted.
Require Import ThieleMachineVerification.ObservationInterface.

(** =========================================================================
    LOCALITY CONSTRAINT
    ========================================================================= *)

(** Partition modules must be spatially local *)
Definition spatial_locality (p : Partition) : Prop :=
  forall m1 m2,
    In m1 p.(modules) ->
    In m2 p.(modules) ->
    m1 <> m2 ->
    (* Disjoint regions - no overlapping spatial support *)
    forall x, In x (snd m1) -> ~ In x (snd m2).

(** =========================================================================
    CAUSALITY CONSTRAINT
    ========================================================================= *)

(** No superluminal influence: module updates cannot affect distant modules
    within a lightcone violation *)
Definition causal_evolution (s s' : ThieleState) : Prop :=
  (* Observable causal constraint at this layer: causal evolution cannot
     arbitrarily change the observable partition signature. *)
  partition_signature s.(partition) = partition_signature s'.(partition).

(** =========================================================================
    UNITARITY / REVERSIBILITY CONSTRAINT
    ========================================================================= *)

(** Information-preserving evolution: blind operations are reversible *)
Definition unitary_evolution (instr : ThieleInstr) : Prop :=
  match instr with
  | EMIT _ => False        (* EMIT is irreversible (measurement) *)
  | HALT => False          (* HALT is irreversible *)
  | PNEW _ _ => True       (* Reversible: can PMERGE *)
  | PSPLIT _ _ _ => True   (* Reversible: can PMERGE *)
  | PMERGE _ _ _ => True   (* Reversible: can PSPLIT *)
  | PDISCOVER _ _ => False (* Sighted operation: information gain *)
  end.

(** =========================================================================
    ENERGY CONSTRAINT (μ as energy)
    ========================================================================= *)

(** Physical evolution conserves or increases μ (no perpetual motion) *)
Definition energy_conservation (s s' : ThieleState) : Prop :=
  s'.(ledger).(mu_total) >= s.(ledger).(mu_total).

(** =========================================================================
    ADMISSIBILITY PREDICATE
    ========================================================================= *)

(** A single instruction is admissible if it satisfies physical constraints *)
Definition instr_admissible (s : ThieleState) (instr : ThieleInstr) (s' : ThieleState) : Prop :=
  spatial_locality s'.(partition) /\
  causal_evolution s s' /\
  energy_conservation s s'.

(** A trace is admissible if every step is admissible *)
Definition trace_has_discover (prog : ThieleProg) : Prop :=
  exists (m : ModuleId) (cost : nat), In (PDISCOVER m cost) prog.

Definition trace_admissible (s : ThieleState) (prog : ThieleProg) : Prop :=
  spatial_locality s.(partition) /\
  (BlindSighted.is_blind_program prog = true \/ trace_has_discover prog).

(** =========================================================================
    ADMISSIBLE SUBSET THEOREMS
    =========================================================================*)

(** Blind programs are always admissible (Turing-complete subset) *)
Theorem blind_programs_admissible : forall s prog,
  spatial_locality s.(partition) ->
  BlindSighted.is_blind_program prog = true ->
  trace_admissible s prog.
Proof.
  intros s prog Hloc Hblind.
  unfold trace_admissible.
  split.
  - exact Hloc.
  - left. exact Hblind.
Qed.

(** =========================================================================
    PHYSICAL LAWS AS THEOREMS
    ========================================================================= *)

(** No-signaling follows from admissibility *)
Theorem admissible_implies_no_signaling : forall s prog,
  trace_admissible s prog ->
  spatial_locality s.(partition).
Proof.
  intros s prog Hadm.
  unfold trace_admissible in Hadm.
  tauto.
Qed.

(** Unitarity of blind evolution *)
Theorem blind_evolution_unitary : forall s prog,
  BlindSighted.is_blind_program prog = true ->
  trace_admissible s prog ->
  BlindSighted.is_blind_program prog = true.
Proof.
  intros s prog Hblind _. exact Hblind.
Qed.

(** =========================================================================
    SIGHTED vs BLIND ADMISSIBILITY
    ========================================================================= *)

(** Sighted operations (PDISCOVER) violate unitarity but preserve causality *)
Theorem pdiscover_breaks_unitarity : forall m cost,
  ~ unitary_evolution (PDISCOVER m cost).
Proof.
  intros m cost.
  unfold unitary_evolution.
  intro Hcontra.
  exact Hcontra.
Qed.

(** But PDISCOVER is still admissible (information gain is physical) *)
Theorem pdiscover_admissible : forall (s : ThieleState) (m : ModuleId * Region) (cost : Z),
  spatial_locality s.(partition) ->
  trace_admissible s [PDISCOVER (fst m) (Z.to_nat cost)].
Proof.
  intros s m cost Hloc.
  unfold trace_admissible.
  split.
  - exact Hloc.
  - right.
    unfold trace_has_discover.
    exists (fst m), (Z.to_nat cost).
    simpl. left. reflexivity.
Qed.

(** =========================================================================
    FALSIFIABILITY
    ========================================================================= *)

(** PREDICTION: Any physical experiment satisfying these admissibility
    constraints must exhibit:
    
    1. No superluminal signaling (from causal_evolution)
    2. Energy conservation (from energy_conservation)  
    3. Spatial locality (from spatial_locality)
    
    EXPERIMENTAL TEST: Violation of any constraint → theory refuted
    *)

(** =========================================================================
    SUMMARY
    ========================================================================= *)

(** This module provides:
    
    1. spatial_locality: modules are spatially disjoint
    2. causal_evolution: no superluminal influence
    3. energy_conservation: μ is monotone increasing
    4. instr_admissible: single-step physical constraint
    5. trace_admissible: full trace satisfies physics
    6. Proven: blind programs are always admissible (TM ⊂ Physics)
    
    Next: Symmetry.v shows which transformations preserve admissibility
    *)
