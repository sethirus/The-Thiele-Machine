From Coq Require Import List Arith.PeanoNat Lia.
Import ListNotations.

Require Import VMState.
Require Import VMStep.
Require Import SimulationProof.

(** * Bounded-model µ-ledger conservation *)

(** The virtual machine executes a bounded trace using [run_vm],
    accumulating µ-costs in the [vm_mu] field of the state.  The ledger
    associated to a bounded execution records, for each realised
    instruction, the µ-delta charged by the specification.  This module
    constructs that ledger and proves that every bounded execution
    preserves the conservation law: the µ-accumulator equals the
    initial µ plus the sum of the recorded deltas, and each consecutive
    pair of states differs exactly by the corresponding ledger entry. *)

(** Ledger extraction from bounded executions. *)

Fixpoint ledger_entries (fuel : nat) (trace : list vm_instruction)
  (s : VMState) : list nat :=
  match fuel with
  | 0 => []
  | S fuel' =>
      match nth_error trace s.(vm_pc) with
      | Some instr =>
          instruction_cost instr ::
          ledger_entries fuel' trace (vm_apply s instr)
      | None => []
      end
  end.

Fixpoint bounded_run (fuel : nat) (trace : list vm_instruction)
  (s : VMState) : list VMState :=
  match fuel with
  | 0 => [s]
  | S fuel' =>
      match nth_error trace s.(vm_pc) with
      | Some instr =>
          s :: bounded_run fuel' trace (vm_apply s instr)
      | None => [s]
      end
  end.

Lemma bounded_run_head :
  forall fuel trace s,
    exists rest, bounded_run fuel trace s = s :: rest.
Proof.
  induction fuel as [|fuel IH]; intros trace s; simpl.
  - exists []. reflexivity.
  - destruct (nth_error trace s.(vm_pc)) as [instr|] eqn:Hlookup.
    + exists (bounded_run fuel trace (vm_apply s instr)). reflexivity.
    + exists []. reflexivity.
Qed.

Lemma vm_apply_mu :
  forall s instr,
    (vm_apply s instr).(vm_mu) = s.(vm_mu) + instruction_cost instr.
Proof.
  intros s instr.
  destruct instr; simpl;
    try (destruct (graph_pnew _ _) as [graph' mid] eqn:?; simpl; reflexivity);
    try (destruct (graph_psplit _ _ _ _) as [[[graph' left_id] right_id]|] eqn:?; simpl; reflexivity);
    try (destruct (graph_pmerge _ _ _) as [[graph' merged_id]|] eqn:?; simpl; reflexivity);
    try (destruct cert as [proof | model]; simpl;
         [destruct (check_lrat formula proof) eqn:?; simpl; reflexivity
         |destruct (check_model formula model) eqn:?; simpl; reflexivity]);
    try (destruct (String.eqb _ _) eqn:?; simpl; reflexivity);
    reflexivity.
Qed.

Fixpoint ledger_conserved (states : list VMState) (entries : list nat)
  : Prop :=
  match states, entries with
  | s :: s' :: rest, delta :: entries' =>
      s'.(vm_mu) = s.(vm_mu) + delta /\
      ledger_conserved (s' :: rest) entries'
  | [_], [] => True
  | _, _ => False
  end.

Lemma ledger_conserved_tail :
  forall s states entries,
    ledger_conserved (s :: states) entries ->
    match states, entries with
    | s' :: rest_states, delta :: rest_entries =>
        s'.(vm_mu) = s.(vm_mu) + delta /\
        ledger_conserved (s' :: rest_states) rest_entries
    | [], [] => True
    | _, _ => False
    end.
Proof.
  intros s states entries H.
  destruct states as [|s' rest].
  - destruct entries as [|delta rest_entries]; simpl in *.
    + exact I.
    + now destruct H.
  - destruct entries as [|delta rest_entries]; simpl in *.
    + now destruct H.
    + destruct H as [Hstep Hrest]. split; auto.
Qed.

(** The next lemma isolates the per-instruction conservation law.
    It asserts that any single small-step transition must debit the
    µ-ledger by exactly the instruction's declared cost.  In particular
    a "free" step—one that changes [vm_mu] without the matching ledger
    delta—would violate [ledger_conserved]; therefore it cannot arise
    under the kernel semantics. *)

Theorem vm_step_respects_mu_ledger :
  forall s instr s',
    vm_step s instr s' ->
    ledger_conserved [s; s'] [instruction_cost instr].
Proof.
  intros s instr s' Hstep.
  simpl.
  split.
  - now apply vm_step_mu.
  - exact I.
Qed.

Fixpoint ledger_sum (entries : list nat) : nat :=
  match entries with
  | [] => 0
  | delta :: rest => delta + ledger_sum rest
  end.

(** ** Irreversibility counting

    Landauer's principle links logically irreversible operations to physical
    entropy production.  To expose that connection, we conservatively count
    irreversible bit events per VM instruction and show the µ-ledger lower
    bounds that count for any bounded execution.  The count is deliberately
    minimal—each instruction contributes at most one irreversible bit and only
    when it charges a positive µ-cost—so the ledger bound holds without extra
    semantic assumptions. *)

Definition irreversible_bits (instr : vm_instruction) : nat :=
  if instruction_cost instr =? 0 then 0 else 1.

Lemma irreversible_bits_le_cost :
  forall instr, irreversible_bits instr <= instruction_cost instr.
Proof.
  intros instr. unfold irreversible_bits.
  destruct (instruction_cost instr =? 0) eqn:Hzero; simpl.
  - apply Nat.eqb_eq in Hzero. subst. lia.
  - apply Nat.eqb_neq in Hzero. lia.
Qed.

Fixpoint irreversible_count (fuel : nat) (trace : list vm_instruction)
  (s : VMState) : nat :=
  match fuel with
  | 0 => 0
  | S fuel' =>
      match nth_error trace s.(vm_pc) with
      | Some instr =>
          irreversible_bits instr +
          irreversible_count fuel' trace (vm_apply s instr)
      | None => 0
      end
  end.

Lemma ledger_sum_bounds_irreversible_count :
  forall fuel trace s,
    irreversible_count fuel trace s <= ledger_sum (ledger_entries fuel trace s).
Proof.
  induction fuel as [|fuel IH]; intros trace s; simpl.
  - lia.
  - destruct (nth_error trace s.(vm_pc)) as [instr|] eqn:Hlookup; simpl.
    + specialize (IH trace (vm_apply s instr)).
      pose proof (irreversible_bits_le_cost instr) as Hbound.
      lia.
    + lia.
Qed.

(** The µ-ledger can now be quoted directly as a bound on the irreversible
    bit events in any bounded execution.  Packaging the previous lemma with a
    more public-facing name makes the Landauer link explicit for downstream
    references. *)

Theorem mu_ledger_bounds_irreversible_events :
  forall fuel trace s,
    irreversible_count fuel trace s <= ledger_sum (ledger_entries fuel trace s).
Proof.
  apply ledger_sum_bounds_irreversible_count.
Qed.

  (** Component-wise accumulation for sighted/blind decompositions.
      The function is parameterised by an instruction-to-cost projection,
      allowing downstream theorems to reason about arbitrary partitions of
    [instruction_cost] (e.g. blind search versus sighted certificates). *)

Fixpoint ledger_component_sum (component : vm_instruction -> nat)
  (fuel : nat) (trace : list vm_instruction) (s : VMState) : nat :=
  match fuel with
  | 0 => 0
  | S fuel' =>
      match nth_error trace s.(vm_pc) with
      | Some instr =>
          component instr +
          ledger_component_sum component fuel' trace (vm_apply s instr)
      | None => 0
      end
  end.

(** Final conservation theorem combining both the cumulative and
    per-step statements. *)

Theorem bounded_model_mu_ledger_conservation :
  forall fuel trace s,
    ledger_conserved (bounded_run fuel trace s)
                     (ledger_entries fuel trace s) /\
  (run_vm fuel trace s).(vm_mu) =
    s.(vm_mu) + ledger_sum (ledger_entries fuel trace s).
Proof.
  induction fuel as [|fuel IH]; intros trace s; simpl.
  - split; [exact I | rewrite Nat.add_0_r; reflexivity].
  - destruct (nth_error trace s.(vm_pc)) as [instr|] eqn:Hlookup; simpl.
    + destruct (IH trace (vm_apply s instr)) as [IH_ledger IH_run].
      destruct (bounded_run_head fuel trace (vm_apply s instr)) as [rest Hrun].
      simpl.
      rewrite Hrun in IH_ledger.
      rewrite Hrun.
      split; [split; [apply vm_apply_mu | exact IH_ledger]
            | rewrite IH_run; rewrite vm_apply_mu; lia].
    + split; [exact I | rewrite Nat.add_0_r; reflexivity].
Qed.

Corollary bounded_ledger_conservation :
  forall fuel trace s,
    ledger_conserved (bounded_run fuel trace s)
                     (ledger_entries fuel trace s).
Proof.
  intros fuel trace s.
  apply (proj1 (bounded_model_mu_ledger_conservation fuel trace s)).
Qed.

Corollary run_vm_mu_conservation :
  forall fuel trace s,
    (run_vm fuel trace s).(vm_mu) =
    s.(vm_mu) + ledger_sum (ledger_entries fuel trace s).
Proof.
  intros fuel trace s.
  apply (proj2 (bounded_model_mu_ledger_conservation fuel trace s)).
Qed.

Corollary run_vm_mu_bounds_irreversibility :
  forall fuel trace s,
    s.(vm_mu) + irreversible_count fuel trace s <= (run_vm fuel trace s).(vm_mu).
Proof.
  intros fuel trace s.
  rewrite run_vm_mu_conservation.
  specialize (ledger_sum_bounds_irreversible_count fuel trace s) as Hbound.
  lia.
Qed.

(** Restating the bound as a delta makes it easier to line up with
    physical arguments about entropy production: the µ-ledger increase over
    an execution interval must dominate the number of irreversible bit
    events recorded by the conservative counter. *)

Theorem run_vm_irreversibility_gap :
  forall fuel trace s,
    irreversible_count fuel trace s <=
      (run_vm fuel trace s).(vm_mu) - s.(vm_mu).
Proof.
  intros fuel trace s.
  rewrite run_vm_mu_conservation.
  specialize (ledger_sum_bounds_irreversible_count fuel trace s) as Hbound.
  lia.
Qed.

(** A quotable alias so downstream developments can refer to the same bound
    without unpacking the µ-delta notation.  This is the flagship lemma for
    mapping µ-ledger growth to a lower bound on logically irreversible bit
    events in a bounded VM execution. *)
Theorem vm_irreversible_bits_lower_bound :
  forall fuel trace s,
    irreversible_count fuel trace s <=
      (run_vm fuel trace s).(vm_mu) - s.(vm_mu).
Proof.
  apply run_vm_irreversibility_gap.
Qed.

Corollary bounded_prefix_mu_balance :
  forall fuel trace s k,
    k <= fuel ->
    (run_vm k trace s).(vm_mu) =
      s.(vm_mu) + ledger_sum (ledger_entries k trace s).
Proof.
  intros fuel trace s k Hle.
  apply run_vm_mu_conservation.
Qed.

(** ** Multi-step µ-monotonicity

    The µ-accumulator never decreases during execution. This follows from
    the fact that [instruction_cost] is always non-negative, ensuring that
    each step either preserves or increases [vm_mu]. *)

Theorem vm_mu_monotonic_single_step :
  forall s instr,
    s.(vm_mu) <= (vm_apply s instr).(vm_mu).
Proof.
  intros s instr.
  rewrite vm_apply_mu.
  lia.
Qed.

Theorem run_vm_mu_monotonic :
  forall fuel trace s,
    s.(vm_mu) <= (run_vm fuel trace s).(vm_mu).
Proof.
  induction fuel as [|fuel IH]; intros trace s; simpl.
  - lia.
  - destruct (nth_error trace s.(vm_pc)) as [instr|] eqn:Hlookup.
    + specialize (IH trace (vm_apply s instr)).
      assert (s.(vm_mu) <= (vm_apply s instr).(vm_mu)) as Hstep.
      { apply vm_mu_monotonic_single_step. }
      lia.
    + lia.
Qed.

(** Extended multi-step monotonicity theorems: The µ-accumulator is preserved
    across execution prefixes and compositional execution phases. *)

Theorem run_vm_mu_monotonic_prefix :
  forall k1 k2 trace s,
    k1 <= k2 ->
    (run_vm k1 trace s).(vm_mu) <= (run_vm k2 trace s).(vm_mu).
Proof.
  intros k1. induction k1 as [|k1 IHk1]; intros k2 trace s Hle.
  - simpl. apply run_vm_mu_monotonic.
  - destruct k2 as [|k2].
    + lia.
    + simpl run_vm.
      destruct (nth_error trace s.(vm_pc)) as [instr|] eqn:Hlookup.
      * apply (IHk1 k2 trace (vm_apply s instr)). lia.
      * simpl. lia.
Qed.

Theorem run_vm_mu_monotonic_composition :
  forall m n trace s,
    s.(vm_mu) <= (run_vm m trace s).(vm_mu) /\
    (run_vm m trace s).(vm_mu) <= (run_vm (m + n) trace s).(vm_mu).
Proof.
  intros m n trace s.
  split.
  - (* First part: s.(vm_mu) <= (run_vm m trace s).(vm_mu) *)
    apply run_vm_mu_monotonic.
  - (* Second part: (run_vm m trace s).(vm_mu) <= (run_vm (m + n) trace s).(vm_mu) *)
    (* Note: run_vm (m + n) = run_vm n (run_vm m s) by the definition of run_vm *)
    assert (forall k1 k2, k1 <= k1 + k2) as Hle by lia.
    apply (run_vm_mu_monotonic_prefix m (m + n) trace s).
    lia.
Qed.

(** We now generalise the conservation statement by splitting the
    instruction cost into complementary components.  This allows the
    kernel development to project the ledger onto semantics such as
    “blind” search work versus “sighted” certificate validation. *)

Section MuDecomposition.

Variable mu_blind_component mu_sighted_component : vm_instruction -> nat.
Variable mu_component_split : forall instr,
  instruction_cost instr =
    mu_blind_component instr + mu_sighted_component instr.

Lemma ledger_sum_component_decompose :
  forall fuel trace s,
    ledger_sum (ledger_entries fuel trace s) =
      ledger_component_sum mu_blind_component fuel trace s +
      ledger_component_sum mu_sighted_component fuel trace s.
Proof.
  induction fuel as [|fuel IH]; intros trace s; simpl.
  - reflexivity.
  - destruct (nth_error trace s.(vm_pc)) as [instr|] eqn:Hlookup.
    + simpl.
      rewrite mu_component_split.
      simpl.
      specialize (IH trace (vm_apply s instr)).
      rewrite IH.
      lia.
    + reflexivity.
Qed.

Theorem bounded_run_mu_decomposition :
  forall fuel trace s,
    (run_vm fuel trace s).(vm_mu) =
      s.(vm_mu) +
      ledger_component_sum mu_blind_component fuel trace s +
      ledger_component_sum mu_sighted_component fuel trace s.
Proof.
  intros fuel trace s.
  destruct (bounded_model_mu_ledger_conservation fuel trace s)
    as [_ Hmu].
  rewrite Hmu.
  rewrite ledger_sum_component_decompose.
  lia.
Qed.

Corollary bounded_run_blind_component_le_total :
  forall fuel trace s,
    s.(vm_mu) + ledger_component_sum mu_blind_component fuel trace s <=
    (run_vm fuel trace s).(vm_mu).
Proof.
  intros fuel trace s.
  rewrite bounded_run_mu_decomposition.
  remember (ledger_component_sum mu_blind_component fuel trace s) as blind_sum.
  remember (ledger_component_sum mu_sighted_component fuel trace s) as sighted_sum.
  lia.
Qed.

Corollary bounded_run_sighted_component_le_total :
  forall fuel trace s,
    s.(vm_mu) + ledger_component_sum mu_sighted_component fuel trace s <=
    (run_vm fuel trace s).(vm_mu).
Proof.
  intros fuel trace s.
  rewrite bounded_run_mu_decomposition.
  remember (ledger_component_sum mu_blind_component fuel trace s) as blind_sum.
  remember (ledger_component_sum mu_sighted_component fuel trace s) as sighted_sum.
  lia.
Qed.

End MuDecomposition.

(** Bridging the prophecy seal and ledger tail.
    The Python experiment derives the gestalt certificate by combining the
    pre-declared seal with the final ledger digest.  The following abstract
    model captures that construction and proves that the gestalt certificate is
    definitionally identical to the computed isomorphism.  The "hash"
    combinator remains uninterpreted here—the property is purely structural and
    does not depend on cryptographic specifics. *)

Section GestaltIsomorphism.

  Variable Hash : Type.
  Variable combine : Hash -> Hash -> Hash.
  Variable default : Hash.

  Definition final_digest (ledger : list Hash) : Hash :=
    match ledger with
    | [] => default
    | _ => List.last ledger default
    end.

  Definition gestalt_certificate (seal : Hash) (ledger : list Hash) : Hash :=
    combine seal (final_digest ledger).

  Definition computed_isomorphism (seal : Hash) (ledger : list Hash) : Hash :=
    combine seal (final_digest ledger).

  Lemma gestalt_matches_isomorphism :
    forall seal ledger,
      gestalt_certificate seal ledger = computed_isomorphism seal ledger.
  Proof.
    intros seal ledger. unfold gestalt_certificate, computed_isomorphism.
    reflexivity.
  Qed.

End GestaltIsomorphism.
