(*
 * ThieleProc: packaging Thiele programs as a process category.
 *
 * This module establishes the first milestone of the geometric
 * unification roadmap: show that Thiele programs with sequential
 * composition form a category.  Objects describe partition interfaces
 * (number of Π-components); morphisms are programs whose receipts run on
 * those interfaces.  Composition is program concatenation and identities
 * are empty programs.  Beyond the category structure we expose helper
 * lemmas about the receipt traces generated by composed programs so later
 * milestones (tensor structure, functors) can reuse them directly.
 *)

From Coq Require Import List Arith.
From ThieleMachine Require Import ThieleMachine.
Import ListNotations.

Set Implicit Arguments.

(* ------------------------------------------------------------------ *)
(* Interfaces *)
(* ------------------------------------------------------------------ *)

Record Interface := {
  iface_partitions : nat;
}.

Definition unit_interface : Interface := {| iface_partitions := 0 |}.

(* Tensor on objects will later become addition on partition counts; we
   introduce the operation now to document the intended geometry even
   though we only need the plain category structure for this milestone. *)
Definition tensor_interface (A B : Interface) : Interface :=
  {| iface_partitions := A.(iface_partitions) + B.(iface_partitions) |}.

(* ------------------------------------------------------------------ *)
(* Programs and sequential composition *)
(* ------------------------------------------------------------------ *)

Definition empty_prog : Prog := {| code := [] |}.

Definition seq_prog (P Q : Prog) : Prog :=
  {| code := P.(code) ++ Q.(code) |}.

Lemma seq_prog_nil_l : forall P, seq_prog empty_prog P = P.
Proof.
  intros [code]. simpl. reflexivity.
Qed.

Lemma seq_prog_nil_r : forall P, seq_prog P empty_prog = P.
Proof.
  intros [instrs]. simpl. apply (f_equal Build_Prog).
  rewrite List.app_nil_r. reflexivity.
Qed.

Lemma seq_prog_assoc : forall P Q R,
  seq_prog (seq_prog P Q) R = seq_prog P (seq_prog Q R).
Proof.
  intros [codeP] [codeQ] [codeR]. simpl.
  apply (f_equal Build_Prog).
  change ((codeP ++ codeQ) ++ codeR = codeP ++ (codeQ ++ codeR)).
  rewrite List.app_assoc. reflexivity.
Qed.

(* ------------------------------------------------------------------ *)
(* Executing programs and observing receipts *)
(* ------------------------------------------------------------------ *)

Definition run_closed (P : Prog) : State * list StepObs :=
  ({| pc := length P.(code) |}, map obs_of_instr P.(code)).

Lemma run_closed_empty :
  run_closed empty_prog = ({| pc := 0 |}, []).
Proof.
  unfold run_closed, empty_prog. simpl. reflexivity.
Qed.

Lemma run_closed_pc : forall P,
  (fst (run_closed P)).(pc) = length P.(code).
Proof.
  intro P. unfold run_closed. simpl. reflexivity.
Qed.


Definition closed_state : State := {| pc := 0 |}.

Fixpoint closed_trace (pc : nat) (instrs : list Instr) : list (State * StepObs) :=
  match instrs with
  | [] => []
  | instr :: tl =>
      ({| pc := S pc |}, obs_of_instr instr) :: closed_trace (S pc) tl
  end.

Definition trace_of_prog (P : Prog) : list (State * StepObs) :=
  closed_trace 0 P.(code).

Fixpoint final_state (s : State) (trace : list (State * StepObs)) : State :=
  match trace with
  | [] => s
  | (s', _) :: tl => final_state s' tl
  end.

Lemma skipn_cons_inv : forall (A : Type) (xs : list A) k a tl,
  skipn k xs = a :: tl ->
  skipn (S k) xs = tl.
Proof.
  intros A xs k. revert xs.
  induction k as [|k IH]; intros xs a tl Hskip.
  - destruct xs as [|x xs]; simpl in Hskip; inversion Hskip; reflexivity.
  - destruct xs as [|x xs]; simpl in Hskip; try discriminate.
    apply IH in Hskip. exact Hskip.
Qed.

Lemma skipn_nth_error : forall (A : Type) (xs : list A) k a tl,
  skipn k xs = a :: tl ->
  nth_error xs k = Some a.
Proof.
  intros A xs k. revert xs.
  induction k as [|k IH]; intros xs a tl Hskip; simpl in *.
  - destruct xs as [|x xs]; inversion Hskip; reflexivity.
  - destruct xs as [|x xs]; simpl in Hskip; try discriminate.
    apply IH in Hskip. exact Hskip.
Qed.

Lemma skipn_succ_suffix : forall (A : Type) (xs : list A) k a tl,
  skipn k xs = a :: tl ->
  skipn (S k) xs = tl.
Proof.
  intros A xs k a tl Hskip.
  apply skipn_cons_inv with (xs:=xs) (a:=a); assumption.
Qed.

Lemma closed_trace_exec_aux : forall P pc suffix,
  skipn pc P.(code) = suffix ->
  Exec P {| pc := pc |} (closed_trace pc suffix).
Proof.
  intros P pc suffix Hskip.
  revert pc Hskip.
  induction suffix as [|instr tl IH]; intros pc Hskip; simpl.
  - constructor.
  - assert (Hnth : nth_error P.(code) pc = Some instr).
    { apply skipn_nth_error with (tl:=tl) in Hskip. exact Hskip. }
    econstructor.
    + apply step_exec. exact Hnth.
    + apply IH. apply skipn_succ_suffix with (a:=instr). exact Hskip.
Qed.

Lemma closed_trace_exec : forall P,
  Exec P closed_state (trace_of_prog P).
Proof.
  intro P. unfold trace_of_prog, closed_state.
  apply closed_trace_exec_aux. simpl. reflexivity.
Qed.
(* Observational equivalence: closed runs produce the same receipts. *)
Definition obs_equiv (P Q : Prog) : Prop :=
  snd (run_closed P) = snd (run_closed Q).

Lemma obs_equiv_refl : forall P, obs_equiv P P.
Proof. intro P. reflexivity. Qed.

Lemma obs_equiv_sym : forall P Q, obs_equiv P Q -> obs_equiv Q P.
Proof. intros P Q H. symmetry. exact H. Qed.

Lemma obs_equiv_trans : forall P Q R,
  obs_equiv P Q -> obs_equiv Q R -> obs_equiv P R.
Proof. intros P Q R HPQ HQR. etransitivity; eauto. Qed.

Lemma run_closed_obs_seq : forall P Q,
  snd (run_closed (seq_prog P Q)) = snd (run_closed P) ++ snd (run_closed Q).
Proof.
  intros [codeP] [codeQ]; simpl. rewrite map_app. reflexivity.
Qed.

Lemma obs_equiv_compose : forall P P' Q Q',
  obs_equiv P P' -> obs_equiv Q Q' ->
  obs_equiv (seq_prog P Q) (seq_prog P' Q').
Proof.
  intros P P' Q Q' HP HQ.
  unfold obs_equiv in *.
  rewrite !run_closed_obs_seq, HP, HQ. reflexivity.
Qed.

Lemma obs_equiv_id_l : forall P,
  obs_equiv (seq_prog empty_prog P) P.
Proof.
  intro P. unfold obs_equiv.
  rewrite run_closed_obs_seq, run_closed_empty. simpl. reflexivity.
Qed.

Lemma obs_equiv_id_r : forall P,
  obs_equiv (seq_prog P empty_prog) P.
Proof.
  intro P. unfold obs_equiv.
  rewrite run_closed_obs_seq, run_closed_empty.
  simpl. rewrite app_nil_r. reflexivity.
Qed.

(* ------------------------------------------------------------------ *)
(* Categorical packaging *)
(* ------------------------------------------------------------------ *)

Record Category := {
  Obj : Type;
  Hom : Obj -> Obj -> Type;
  id  : forall {A}, Hom A A;
  comp : forall {A B C}, Hom B C -> Hom A B -> Hom A C;
  comp_assoc : forall A B C D (h : Hom C D) (g : Hom B C) (f : Hom A B),
      comp h (comp g f) = comp (comp h g) f;
  comp_id_left : forall A B (f : Hom A B), comp (@id B) f = f;
  comp_id_right : forall A B (f : Hom A B), comp f (@id A) = f
}.

Definition ThieleProc : Category :=
  {| Obj := Interface;
     Hom _ _ := Prog;
     id _ := empty_prog;
     comp _ _ _ g f := seq_prog f g;
     comp_assoc _ _ _ _ h g f := seq_prog_assoc f g h;
     comp_id_left _ _ f := seq_prog_nil_r f;
     comp_id_right _ _ f := seq_prog_nil_l f |}.

(* ------------------------------------------------------------------ *)
(* Interface helpers for upcoming tensor proofs *)
(* ------------------------------------------------------------------ *)

Lemma iface_tensor_partitions : forall A B,
  (tensor_interface A B).(iface_partitions) =
  A.(iface_partitions) + B.(iface_partitions).
Proof.
  intros A B. reflexivity.
Qed.

Lemma run_closed_tensor_pc : forall P Q,
  (fst (run_closed (seq_prog P Q))).(pc) =
    (fst (run_closed P)).(pc) + (fst (run_closed Q)).(pc).
Proof.
  intros P Q. unfold run_closed, seq_prog. simpl. rewrite app_length. reflexivity.
Qed.

(* The lemmas above give the concrete footholds required by the remaining
   milestones: tensor structure (running programs in parallel) and
   embeddings from logic/computation/physics.  Later files will build on
   `ThieleProc` rather than re-developing sequential reasoning. *)
