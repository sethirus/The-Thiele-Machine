// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// Copyright 2025 Devon Thiele
// See the LICENSE file in the repository root for full terms.

// ============================================================================
// Thiele CPU Python Execution Engine (PEE)
// ============================================================================

module pee (
    input wire clk,
    input wire rst_n,

    // CPU interface
    input wire py_req,
    input wire [31:0] py_code_addr,
    output wire py_ack,
    output wire [31:0] py_result,

    // External Python interface
    output wire python_req,
    output wire [31:0] python_code_addr,
    input wire python_ack,
    input wire [31:0] python_result,
    input wire python_error,

    // Symbolic execution interface
    output wire symbolic_req,
    output wire [31:0] symbolic_vars,
    input wire symbolic_ack,
    input wire [31:0] symbolic_assignment,

    // Status
    output wire [31:0] pee_status,
    output wire pee_error
);

// ============================================================================
// PARAMETERS AND STATES
// ============================================================================

localparam STATE_IDLE = 3'h0;
localparam STATE_LOAD_CODE = 3'h1;
localparam STATE_EXECUTE = 3'h2;
localparam STATE_SYMBOLIC = 3'h3;
localparam STATE_WAIT_RESULT = 3'h4;
localparam STATE_COMPLETE = 3'h5;

// Error codes
localparam ERR_NONE = 32'h0;
localparam ERR_TIMEOUT = 32'h4001;
localparam ERR_PYTHON_ERROR = 32'h4002;
localparam ERR_SYMBOLIC_FAIL = 32'h4003;

// ============================================================================
// INTERNAL REGISTERS
// ============================================================================

reg [2:0] state;
reg [31:0] current_code_addr;
reg [31:0] execution_result;
reg ack_pending;
reg [15:0] timeout_counter;
reg [31:0] error_code;

// Symbolic execution state
reg [31:0] symbolic_var_count;
reg [31:0] symbolic_domain_size;
reg symbolic_mode;

// Execution statistics
reg [31:0] execution_count;
reg [31:0] symbolic_count;
reg [31:0] error_count;

// ============================================================================
// CODE ANALYSIS LOGIC
// ============================================================================

wire is_symbolic_code;
wire [31:0] var_count;
wire [31:0] domain_size;

// Simple code analysis (would be more sophisticated in real implementation)
assign is_symbolic_code = (py_code_addr[31:28] == 4'hA); // Marker for symbolic code
assign var_count = py_code_addr[27:24]; // Encoded variable count
assign domain_size = py_code_addr[23:20]; // Encoded domain size

// ============================================================================
// STATE MACHINE
// ============================================================================

always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        state <= STATE_IDLE;
        ack_pending <= 1'b0;
        timeout_counter <= 16'h0;
        error_code <= ERR_NONE;
        execution_result <= 32'h0;
        symbolic_var_count <= 32'h0;
        symbolic_domain_size <= 32'h0;
        symbolic_mode <= 1'b0;
        execution_count <= 32'h0;
        symbolic_count <= 32'h0;
        error_count <= 32'h0;
    end else begin
        case (state)
            STATE_IDLE: begin
                if (py_req && !ack_pending) begin
                    current_code_addr <= py_code_addr;
                    timeout_counter <= 16'hFFFF; // ~1ms timeout
                    error_code <= ERR_NONE;

                    if (is_symbolic_code) begin
                        state <= STATE_SYMBOLIC;
                        symbolic_mode <= 1'b1;
                        symbolic_var_count <= var_count;
                        symbolic_domain_size <= domain_size;
                    end else begin
                        state <= STATE_LOAD_CODE;
                        symbolic_mode <= 1'b0;
                    end
                end
            end

            STATE_LOAD_CODE: begin
                state <= STATE_EXECUTE;
            end

            STATE_EXECUTE: begin
                state <= STATE_WAIT_RESULT;
            end

            STATE_SYMBOLIC: begin
                state <= STATE_WAIT_RESULT;
            end

            STATE_WAIT_RESULT: begin
                timeout_counter <= timeout_counter - 1;

                if (symbolic_mode ? symbolic_ack : python_ack) begin
                    if (symbolic_mode) begin
                        execution_result <= symbolic_assignment;
                        symbolic_count <= symbolic_count + 1;
                    end else begin
                        execution_result <= python_result;
                        execution_count <= execution_count + 1;

                        if (python_error) begin
                            error_code <= ERR_PYTHON_ERROR;
                            error_count <= error_count + 1;
                        end
                    end

                    state <= STATE_COMPLETE;
                    ack_pending <= 1'b1;

                end else if (timeout_counter == 0) begin
                    state <= STATE_COMPLETE;
                    error_code <= ERR_TIMEOUT;
                    error_count <= error_count + 1;
                    ack_pending <= 1'b1;
                end
            end

            STATE_COMPLETE: begin
                if (!py_req) begin
                    state <= STATE_IDLE;
                    ack_pending <= 1'b0;
                    symbolic_mode <= 1'b0;
                end
            end

            default: begin
                state <= STATE_IDLE;
            end
        endcase
    end
end

// ============================================================================
// SYMBOLIC EXECUTION LOGIC
// ============================================================================

wire [31:0] total_combinations;
wire [31:0] symbolic_domain_n;
wire [31:0] symbolic_domain_mask;

// Domain size encoding is interpreted as an exponent: domain_n = 2^domain_size.
// This keeps the symbolic assignment generator synthesizable (no variable '%').
assign symbolic_domain_n = (symbolic_domain_size < 32) ? (32'h1 << symbolic_domain_size[4:0]) : 32'h0;
assign symbolic_domain_mask = (symbolic_domain_n == 0) ? 32'h0 : (symbolic_domain_n - 1);
assign total_combinations = symbolic_var_count * symbolic_domain_n;

// Simple symbolic solver (brute force for demonstration)
reg [31:0] current_try;
reg [31:0] assignment;

always @(posedge clk) begin
    if (state == STATE_SYMBOLIC) begin
        // Generate next assignment to try
        current_try <= current_try + 1;
        assignment <= current_try & symbolic_domain_mask;
    end else begin
        current_try <= 32'h0;
        assignment <= 32'h0;
    end
end

// ============================================================================
// OUTPUT ASSIGNMENTS
// ============================================================================

assign python_req = (state == STATE_EXECUTE);
assign python_code_addr = current_code_addr;
assign symbolic_req = (state == STATE_SYMBOLIC);
assign symbolic_vars = {symbolic_var_count[15:0], symbolic_domain_size[15:0]};
assign py_ack = ack_pending;
assign py_result = execution_result;
assign pee_status = {execution_count[15:0], symbolic_count[15:0]};
assign pee_error = (error_code != ERR_NONE);

endmodule