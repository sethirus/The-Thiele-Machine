(* ================================================================= *)
(* Thiele Machine Concrete Pack - Module Packaging *)
(* ================================================================= *)

(* This file depends on ThieleMachineUniv.v which has module issues.
   The MAIN WORKING IMPLEMENTATION is in ThieleMachineConcrete.v.
   
   For the verified implementation, see:
   - coq/thielemachine/coqproofs/ThieleMachineConcrete.v (WORKING)
   - coq/thielemachine/coqproofs/Subsumption.v (main theorems, PROVEN)
   - docs/FIXED_FILES_SUMMARY.md (compilation status) *)
