(** =========================================================================
    CORE SEMANTICS - Canonical Formal Specification
    =========================================================================
    
    This module provides the canonical, self-contained formal semantics
    for the Thiele Machine as specified in docs/MODEL_SPEC.md (A1.2).
    
    This file implements Task A1.3 from the Research Program Master Plan:
    - Complete formal state space S
    - Transition system (step function)
    - Multi-step execution (run function)
    - μ-cost accounting (μ-update function)
    
    DESIGN PRINCIPLES:
    1. Self-contained: No external dependencies except Coq stdlib
    2. Executable: All definitions computable
    3. Verifiable: All claims proven with Qed
    4. Aligned: Matches Python VM (thielecpu/) and Verilog (hardware/)
    
    STATUS: Task A1.3 (Create Formal Semantics) - COMPLETE
    NEXT: Task A1.4 (Prove Core Invariants)
    
    =========================================================================
    REFERENCES
    =========================================================================
    
    [MODEL_SPEC] docs/MODEL_SPEC.md - Canonical model specification
    [PYTHON_VM] thielecpu/vm.py - Reference implementation
    [VERILOG] thielecpu/hardware/thiele_cpu.v - Hardware implementation
    [BLIND_SIGHTED] BlindSighted.v - Blind/Sighted separation
    [THIELE_MACHINE] ThieleMachine.v - Abstract machine interface
    
    ========================================================================= *)

From Coq Require Import List String ZArith Lia Bool Nat.
Require Import ThieleMachine.Hash256.
Import ListNotations.
Open Scope Z_scope.

(** =========================================================================
    SECTION 1: STATE SPACE S
    =========================================================================
    
    The state space S consists of:
    - Variables and their assignments
    - Partitions (modules dividing the state space)
    - μ-ledger (information cost accounting)
    - Program counter and control flow state
    
    ========================================================================= *)

(** Basic types *)
Definition VarId := nat.
Definition ModuleId := nat.
Definition Region := list VarId.

(** Partition: A collection of disjoint modules *)
Record Partition := {
  modules : list (ModuleId * Region);
  next_module_id : ModuleId;
}.

(** Empty partition (initialization) *)
Definition empty_partition : Partition :=
  {| modules := [];
     next_module_id := 0%nat |}.

(** Trivial partition: all variables in one module *)
Definition trivial_partition (vars : Region) : Partition :=
  {| modules := [(0%nat, vars)];
     next_module_id := 1%nat |}.

(** μ-Ledger: Tracks information cost *)
Record MuLedger := {
  mu_operational : Z;    (* Cost of computation steps *)
  mu_information : Z;    (* Cost of information revelation *)
  mu_total : Z;          (* Total cost = operational + information *)
}.

(** Zero ledger (initial state) *)
Definition zero_mu : MuLedger :=
  {| mu_operational := 0;
     mu_information := 0;
     mu_total := 0 |}.

(** Add operational cost *)
Definition add_mu_operational (l : MuLedger) (delta : Z) : MuLedger :=
  {| mu_operational := l.(mu_operational) + delta;
     mu_information := l.(mu_information);
     mu_total := l.(mu_total) + delta |}.

(** Add information cost *)
Definition add_mu_information (l : MuLedger) (delta : Z) : MuLedger :=
  {| mu_operational := l.(mu_operational);
     mu_information := l.(mu_information) + delta;
     mu_total := l.(mu_total) + delta |}.

(** Instruction set - defined before State to avoid forward reference *)
Inductive Instruction : Type :=
  | PNEW : Region -> Instruction              (* 0x00: Create module *)
  | PSPLIT : ModuleId -> Instruction          (* 0x01: Split module *)
  | PMERGE : ModuleId -> ModuleId -> Instruction  (* 0x02: Merge modules *)
  | LASSERT : Instruction                     (* 0x03: Logical assertion *)
  | LJOIN : Instruction                       (* 0x04: Logical join *)
  | MDLACC : ModuleId -> Instruction          (* 0x05: Accumulate MDL *)
  | PDISCOVER : Instruction                   (* 0x06: Discover partition *)
  | XFER : Instruction                        (* 0x07: Transfer *)
  | PYEXEC : Instruction                      (* 0x08: Python execution *)
  | XOR_LOAD : Instruction                    (* 0x0A: XOR load *)
  | XOR_ADD : Instruction                     (* 0x0B: XOR add *)
  | XOR_SWAP : Instruction                    (* 0x0C: XOR swap *)
  | XOR_RANK : Instruction                    (* 0x0D: XOR rank *)
  | EMIT : nat -> Instruction                 (* 0x0E: Emit result *)
  | ORACLE_HALTS : Instruction                (* 0x0F: Oracle halting *)
  | HALT : Instruction.                       (* 0xFF: Halt *)

(** Program: List of instructions *)
Definition Program := list Instruction.

(** Complete Thiele Machine State *)
Record State := {
  partition : Partition;    (* Current partition structure *)
  mu_ledger : MuLedger;     (* μ-cost accumulator *)
  pc : nat;                 (* Program counter *)
  halted : bool;            (* Halting flag *)
  result : option nat;      (* Final result *)
  program : Program;        (* Program being executed *)
}.

(** Initial state *)
Definition initial_state (vars : Region) (prog : Program) : State :=
  {| partition := trivial_partition vars;
     mu_ledger := zero_mu;
     pc := 0;
     halted := false;
     result := None;
     program := prog |}.

(** =========================================================================
    SECTION 1.5: CRYPTOGRAPHIC RECEIPTS INFRASTRUCTURE
    =========================================================================
    
    To prevent receipt forgery, we add cryptographic binding via state hashes.
    Each execution step creates a cryptographic commitment to the complete state.
    These commitments form a hash chain that binds the receipt to the actual
    execution path.
    
    KEY PROPERTY: By collision resistance of the hash function, forging a valid
    receipt requires finding states that hash to the committed values and follow
    valid transition rules - computationally equivalent to honest execution.
    
    ========================================================================= *)

(** State hash: 256-bit cryptographic commitment to state 
    Represented as list of 256 booleans (bits)
    
    BIT ORDERING: Big-endian (MSB first)
    - Position 0 = most significant bit
    - Position 255 = least significant bit
    
    CANONICAL ENCODING: States are serialized deterministically as:
    1. Partition: sorted list of (module_id, sorted_variables)
    2. μ-ledger: (mu_operational, mu_information, mu_total) as big-endian Z
    3. PC: nat as big-endian
    4. Halted: 0 or 1
    5. Result: None = 0x00, Some(n) = 0x01 || n
    6. Program: SHA-256 hash of program (not full program)
    
    This encoding MUST match Python hash_snapshot() and Verilog state_hasher
    for cross-layer isomorphism.
*)
Definition StateHash := list bool.

(** Hash function: State -> 256-bit commitment.

    This is an *executable* deterministic hash inside Coq (no Parameters/Axioms).
    It is NOT a cryptographic hash. If you need cryptographic guarantees, keep
    them as external claims and validate SHA-256 alignment in the Python/Verilog
    pipeline.
*)

Definition bool_to_Z (b : bool) : Z := if b then 1 else 0.

Fixpoint encode_region (r : Region) : list Z :=
  match r with
  | [] => []
  | x :: xs => Z.of_nat x :: encode_region xs
  end.

Fixpoint encode_modules (ms : list (ModuleId * Region)) : list Z :=
  match ms with
  | [] => []
  | (mid, r) :: ms' =>
      Z.of_nat mid :: Z.of_nat (List.length r) :: encode_region r ++ encode_modules ms'
  end.

Definition encode_partition (p : Partition) : list Z :=
  encode_modules p.(modules) ++ [Z.of_nat p.(next_module_id)].

Definition instr_tag (i : Instruction) : Z :=
  match i with
  | PNEW _ => 0
  | PSPLIT _ => 1
  | PMERGE _ _ => 2
  | LASSERT => 3
  | LJOIN => 4
  | MDLACC _ => 5
  | PDISCOVER => 6
  | XFER => 7
  | PYEXEC => 8
  | XOR_LOAD => 10
  | XOR_ADD => 11
  | XOR_SWAP => 12
  | XOR_RANK => 13
  | EMIT _ => 14
  | ORACLE_HALTS => 15
  | HALT => 255
  end.

Definition encode_instruction (i : Instruction) : list Z :=
  match i with
  | PNEW r => [instr_tag i; Z.of_nat (List.length r)] ++ encode_region r
  | PSPLIT m => [instr_tag i; Z.of_nat m]
  | PMERGE m1 m2 => [instr_tag i; Z.of_nat m1; Z.of_nat m2]
  | MDLACC m => [instr_tag i; Z.of_nat m]
  | EMIT n => [instr_tag i; Z.of_nat n]
  | _ => [instr_tag i]
  end.

Fixpoint encode_program (p : Program) : list Z :=
  match p with
  | [] => []
  | i :: ps => encode_instruction i ++ encode_program ps
  end.

Definition encode_state (s : State) : list Z :=
  encode_partition s.(partition)
  ++ [s.(mu_ledger).(mu_operational); s.(mu_ledger).(mu_information); s.(mu_ledger).(mu_total)]
  ++ [Z.of_nat s.(pc); bool_to_Z s.(halted)]
  ++ (match s.(result) with None => [0] | Some n => [1; Z.of_nat n] end)
  ++ [Z.of_nat (List.length s.(program))]
  ++ encode_program s.(program).

Definition hash_state (s : State) : StateHash := Hash256.hash256 (encode_state s).

(** Helper: Compare state hashes for equality
    
    NOTE: This recursive implementation performs 256 comparisons for full hash.
    For actual implementations (Python/Verilog), use optimized equality:
    - Python: h1 == h2 (native string/bytes comparison)
    - Verilog: assign equal = (h1 == h2); (hardware parallel comparison)
    
    The recursive Fixpoint is used here for Coq reasoning and proof simplicity.
*)
Fixpoint hash_eq (h1 h2 : StateHash) : bool :=
  match h1, h2 with
  | [], [] => true
  | b1 :: h1', b2 :: h2' => Bool.eqb b1 b2 && hash_eq h1' h2'
  | _, _ => false
  end.

(** =========================================================================
    SECTION 2: INSTRUCTION SET
    =========================================================================
    
    Core instructions aligned with Python VM and Verilog RTL:
    - PNEW: Create partition module
    - PSPLIT: Split module
    - PMERGE: Merge modules
    - PDISCOVER: Auto-discover partition
    - LASSERT: Logical assertion
    - MDLACC: MDL cost accumulation
    - EMIT: Emit result
    - HALT: Stop execution
    
    Opcode alignment:
    - Python: thielecpu/isa.py
    - Verilog: thielecpu/hardware/thiele_cpu.v (OPCODE_* parameters)
    - Coq: This file
    
    ========================================================================= *)

(** Note: Instruction and Program types defined earlier (before State record) *)

(** =========================================================================
    SECTION 3: TRANSITION SYSTEM (STEP FUNCTION)
    =========================================================================
    
    Small-step operational semantics: step : State -> option State
    
    Each instruction updates:
    1. Partition (for PNEW, PSPLIT, PMERGE, PDISCOVER)
    2. μ-ledger (all instructions incur cost)
    3. Program counter (incremented or halt)
    4. Result (for EMIT)
    
    Returns None if execution cannot proceed (already halted).
    
    ========================================================================= *)

(** Helper: Add a module to partition *)
Definition add_module (p : Partition) (r : Region) : Partition :=
  {| modules := p.(modules) ++ [(p.(next_module_id), r)];
     next_module_id := S p.(next_module_id) |}.

(** Region equality and overlap checks (used to enforce partition validity for PNEW). *)
Fixpoint region_eqb (r1 r2 : Region) : bool :=
  match r1, r2 with
  | [], [] => true
  | x :: xs, y :: ys => Nat.eqb x y && region_eqb xs ys
  | _, _ => false
  end.

Definition region_overlap_b (r1 r2 : Region) : bool :=
  existsb (fun x => existsb (Nat.eqb x) r2) r1.

Lemma region_eqb_refl : forall r, region_eqb r r = true.
Proof.
  induction r as [|x xs IH]; simpl; auto.
  rewrite Nat.eqb_refl. rewrite IH. reflexivity.
Qed.

(** Helper: Find module by ID *)
Fixpoint find_module_in_list (mods : list (ModuleId * Region)) (mid : ModuleId) : option Region :=
  match mods with
  | [] => None
  | (id, r) :: rest =>
      if Nat.eqb id mid then Some r
      else find_module_in_list rest mid
  end.

Definition find_module (p : Partition) (mid : ModuleId) : option Region :=
  find_module_in_list p.(modules) mid.

(** Lemma: find_module_in_list preserves lookups when appending *)
Lemma find_module_in_list_app : forall mods mid new_entry,
  (forall id r, In (id, r) [new_entry] -> id <> mid) ->
  find_module_in_list (mods ++ [new_entry]) mid = find_module_in_list mods mid.
Proof.
  intros mods mid new_entry Hnew.
  induction mods as [| [id r] rest IH].
  - (* Base case: empty list *)
    simpl.
    destruct new_entry as [new_id new_r].
    destruct (Nat.eqb new_id mid) eqn:Heq.
    + (* new_id = mid, contradiction *)
      apply Nat.eqb_eq in Heq.
      exfalso.
      apply (Hnew new_id new_r).
      * simpl. left. reflexivity.
      * assumption.
    + (* new_id <> mid, return None *)
      reflexivity.
  - (* Inductive case *)
    simpl.
    destruct (Nat.eqb id mid) eqn:Heq.
    + (* Found it, return immediately *)
      reflexivity.
    + (* Not found, recurse *)
      apply IH.
Qed.

(** Lemma: add_module preserves existing module lookups *)
Lemma add_module_preserves : forall p r mid,
  (mid < p.(next_module_id))%nat ->
  find_module (add_module p r) mid = find_module p mid.
Proof.
  intros p r mid Hlt.
  unfold add_module, find_module. simpl.
  apply find_module_in_list_app.
  intros id reg Hin.
  simpl in Hin.
  destruct Hin as [Heq | Hfalse].
  - (* The new entry has id = next_module_id *)
    injection Heq as Heq_id Heq_r.
    subst id.
    (* next_module_id > mid by assumption *)
    (* mid < next_module_id means mid <> next_module_id *)
    intros Heq_contra.
    rewrite Heq_contra in Hlt.
    apply Nat.lt_irrefl in Hlt.
    exact Hlt.
  - (* No other entries in the singleton list *)
    contradiction.
Qed.

(** Helper: Split a region into even and odd variables *)
Definition split_region (r : Region) : Region * Region :=
  List.partition Nat.even r.

(** Helper: Remove a module from the list *)
Fixpoint remove_module_from_list (mods : list (ModuleId * Region)) (mid : ModuleId) : list (ModuleId * Region) :=
  match mods with
  | [] => []
  | (id, r) :: rest =>
      if Nat.eqb id mid then rest
      else (id, r) :: remove_module_from_list rest mid
  end.

(** Helper: Update partition for PSPLIT *)
Definition update_partition_split (p : Partition) (mid : ModuleId) : Partition :=
  match find_module p mid with
  | None => p
  | Some r =>
      let (r_even, r_odd) := split_region r in
      let mods' := remove_module_from_list p.(modules) mid in
      let id1 := p.(next_module_id) in
      let id2 := S p.(next_module_id) in
      {| modules := mods' ++ [(id1, r_even); (id2, r_odd)];
         next_module_id := S (S p.(next_module_id)) |}
  end.

(** Helper: Update partition for PMERGE *)
Definition update_partition_merge (p : Partition) (m1 m2 : ModuleId) : Partition :=
  match find_module p m1, find_module p m2 with
  | Some r1, Some r2 =>
      let mods' := remove_module_from_list (remove_module_from_list p.(modules) m1) m2 in
      let new_id := p.(next_module_id) in
      {| modules := mods' ++ [(new_id, r1 ++ r2)];
         next_module_id := S p.(next_module_id) |}
  | _, _ => p
  end.

(** Helper: Boolean disjointness check *)
Definition disjoint_b (r1 r2 : Region) : bool :=
  forallb (fun x => negb (existsb (Nat.eqb x) r2)) r1.

(** Helper: Boolean partition validity check *)
Fixpoint regions_disjoint_b (regions : list Region) : bool :=
  match regions with
  | [] => true
  | r :: rest =>
      (forallb (fun r' => disjoint_b r r') rest) &&
      regions_disjoint_b rest
  end.

Definition partition_valid_b (p : Partition) : bool :=
  regions_disjoint_b (map snd p.(modules)).

(** μ-cost for partition operations (from μ-spec v2.0) *)
Definition mu_pnew_cost : Z := 8.     (* Cost to create module *)
Definition mu_psplit_cost : Z := 16.  (* Cost to split module *)
Definition mu_pmerge_cost : Z := 12.  (* Cost to merge modules *)
Definition mu_pdiscover_cost : Z := 100. (* Cost to discover partition *)
Definition mu_lassert_cost : Z := 20. (* Cost for logical assertion *)
Definition mu_mdlacc_cost : Z := 5.   (* Cost for MDL accumulation *)
Definition mu_emit_cost : Z := 1.     (* Cost to emit result *)

Lemma mu_pnew_cost_nonneg : 0 <= mu_pnew_cost.
Proof. cbv [mu_pnew_cost]. lia. Qed.

Lemma mu_psplit_cost_nonneg : 0 <= mu_psplit_cost.
Proof. cbv [mu_psplit_cost]. lia. Qed.

Lemma mu_pmerge_cost_nonneg : 0 <= mu_pmerge_cost.
Proof. cbv [mu_pmerge_cost]. lia. Qed.

Lemma mu_pdiscover_cost_nonneg : 0 <= mu_pdiscover_cost.
Proof. cbv [mu_pdiscover_cost]. lia. Qed.

Lemma mu_lassert_cost_nonneg : 0 <= mu_lassert_cost.
Proof. cbv [mu_lassert_cost]. lia. Qed.

Lemma mu_mdlacc_cost_nonneg : 0 <= mu_mdlacc_cost.
Proof. cbv [mu_mdlacc_cost]. lia. Qed.

Lemma mu_emit_cost_nonneg : 0 <= mu_emit_cost.
Proof. cbv [mu_emit_cost]. lia. Qed.

Lemma add_mu_operational_mu_total_ge :
  forall (l : MuLedger) (delta : Z),
    0 <= delta ->
    (add_mu_operational l delta).(mu_total) >= l.(mu_total).
Proof.
  intros l delta Hdelta.
  unfold add_mu_operational. simpl.
  lia.
Qed.

Lemma add_mu_information_mu_total_ge :
  forall (l : MuLedger) (delta : Z),
    0 <= delta ->
    (add_mu_information l delta).(mu_total) >= l.(mu_total).
Proof.
  intros l delta Hdelta.
  unfold add_mu_information. simpl.
  lia.
Qed.

(** Single-step execution *)
Definition step (s : State) : option State :=
  if s.(halted) then None  (* Cannot step if halted *)
  else
    match nth_error s.(program) s.(pc) with
    | None => Some {| partition := s.(partition);
                      mu_ledger := s.(mu_ledger);
                      pc := s.(pc);
                      halted := true;
                      result := s.(result);
                      program := s.(program) |}  (* Halt if PC out of bounds *)
    | Some instr =>
        match instr with
        | PNEW r =>
          (* Create new partition module.
             Canonical semantics (per MODEL_SPEC):
             - Deduplicate exact duplicates (no-op, Δμ=0)
             - Reject partial overlaps (halt)
             - Otherwise add disjoint region.
          *)
          let regs := map snd s.(partition).(modules) in
          if existsb (fun r' => region_eqb r r') regs then
            (* Exact duplicate: no-op *)
            Some {| partition := s.(partition);
              mu_ledger := s.(mu_ledger);
              pc := S s.(pc);
              halted := false;
              result := s.(result);
              program := s.(program) |}
          else if existsb (fun r' => negb (disjoint_b r r')) regs then
            (* Partial overlap: halt (preserves validity) *)
            Some {| partition := s.(partition);
              mu_ledger := s.(mu_ledger);
              pc := s.(pc);
              halted := true;
              result := None;
              program := s.(program) |}
          else
            (* New disjoint region: add it and charge μ (only if validity holds). *)
            let p' := add_module s.(partition) r in
            if partition_valid_b p' then
              let mu' := add_mu_operational s.(mu_ledger) mu_pnew_cost in
              Some {| partition := p';
                mu_ledger := mu';
                pc := S s.(pc);
                halted := false;
                result := s.(result);
                program := s.(program) |}
            else
              (* Defensive: refuse to enter an invalid partition state. *)
              Some {| partition := s.(partition);
                mu_ledger := s.(mu_ledger);
                pc := s.(pc);
                halted := true;
                result := None;
                program := s.(program) |}
        
        | PSPLIT mid =>
            (* Split module: Even/Odd split *)
            let p' := update_partition_split s.(partition) mid in
            if partition_valid_b p' then
              let mu' := add_mu_operational s.(mu_ledger) mu_psplit_cost in
              Some {| partition := p';
                mu_ledger := mu';
                pc := S s.(pc);
                halted := false;
                result := s.(result);
                program := s.(program) |}
            else
              (* Defensive: refuse to enter an invalid partition state, but still charge μ for the attempted split. *)
              let mu' := add_mu_operational s.(mu_ledger) mu_psplit_cost in
              Some {| partition := s.(partition);
                mu_ledger := mu';
                pc := s.(pc);
                halted := true;
                result := None;
                program := s.(program) |}
        
        | PMERGE m1 m2 =>
            (* Merge modules *)
            let p' := update_partition_merge s.(partition) m1 m2 in
            if partition_valid_b p' then
              let mu' := add_mu_operational s.(mu_ledger) mu_pmerge_cost in
              Some {| partition := p';
                mu_ledger := mu';
                pc := S s.(pc);
                halted := false;
                result := s.(result);
                program := s.(program) |}
            else
              (* Defensive: refuse to enter an invalid partition state. *)
              Some {| partition := s.(partition);
                mu_ledger := s.(mu_ledger);
                pc := s.(pc);
                halted := true;
                result := None;
                program := s.(program) |}

        | PDISCOVER =>
            (* Auto-discover partition *)
            let mu' := add_mu_information s.(mu_ledger) mu_pdiscover_cost in
            Some {| partition := s.(partition);
                    mu_ledger := mu';
                    pc := S s.(pc);
                    halted := false;
                    result := s.(result);
                    program := s.(program) |}

        | LASSERT =>
            (* Logical assertion: Check partition validity *)
            if partition_valid_b s.(partition) then
              let mu' := add_mu_operational s.(mu_ledger) mu_lassert_cost in
              Some {| partition := s.(partition);
                      mu_ledger := mu';
                      pc := S s.(pc);
                      halted := false;
                      result := s.(result);
                      program := s.(program) |}
            else
              (* Assertion failed: Halt *)
              Some {| partition := s.(partition);
                      mu_ledger := s.(mu_ledger);
                      pc := s.(pc);
                      halted := true;
                      result := None;
                      program := s.(program) |}

        | LJOIN =>
            (* Logical join *)
            let mu' := add_mu_operational s.(mu_ledger) mu_lassert_cost in
            Some {| partition := s.(partition);
                    mu_ledger := mu';
                    pc := S s.(pc);
                    halted := false;
                    result := s.(result);
                    program := s.(program) |}

        | MDLACC mid =>
            (* MDL cost accumulation *)
            let mu' := add_mu_operational s.(mu_ledger) mu_mdlacc_cost in
            Some {| partition := s.(partition);
                    mu_ledger := mu';
                    pc := S s.(pc);
                    halted := false;
                    result := s.(result);
                    program := s.(program) |}

        | XFER =>
            (* Transfer operation *)
            let mu' := add_mu_operational s.(mu_ledger) mu_emit_cost in
            Some {| partition := s.(partition);
                    mu_ledger := mu';
                    pc := S s.(pc);
                    halted := false;
                    result := s.(result);
                    program := s.(program) |}

        | PYEXEC =>
            (* Python execution *)
            let mu' := add_mu_operational s.(mu_ledger) mu_lassert_cost in
            Some {| partition := s.(partition);
                    mu_ledger := mu';
                    pc := S s.(pc);
                    halted := false;
                    result := s.(result);
                    program := s.(program) |}

        | XOR_LOAD =>
            (* XOR load operation *)
            let mu' := add_mu_operational s.(mu_ledger) mu_emit_cost in
            Some {| partition := s.(partition);
                    mu_ledger := mu';
                    pc := S s.(pc);
                    halted := false;
                    result := s.(result);
                    program := s.(program) |}

        | XOR_ADD =>
            (* XOR add operation *)
            let mu' := add_mu_operational s.(mu_ledger) mu_emit_cost in
            Some {| partition := s.(partition);
                    mu_ledger := mu';
                    pc := S s.(pc);
                    halted := false;
                    result := s.(result);
                    program := s.(program) |}

        | XOR_SWAP =>
            (* XOR swap operation *)
            let mu' := add_mu_operational s.(mu_ledger) mu_emit_cost in
            Some {| partition := s.(partition);
                    mu_ledger := mu';
                    pc := S s.(pc);
                    halted := false;
                    result := s.(result);
                    program := s.(program) |}

        | XOR_RANK =>
            (* XOR rank operation *)
            let mu' := add_mu_operational s.(mu_ledger) mu_emit_cost in
            Some {| partition := s.(partition);
                    mu_ledger := mu';
                    pc := S s.(pc);
                    halted := false;
                    result := s.(result);
                    program := s.(program) |}

        | EMIT n =>
            (* Emit result *)
            let mu' := add_mu_operational s.(mu_ledger) mu_emit_cost in
            Some {| partition := s.(partition);
                    mu_ledger := mu';
                    pc := S s.(pc);
                    halted := false;
                    result := Some n;
                    program := s.(program) |}

        | ORACLE_HALTS =>
            (* Oracle halting check *)
            let mu' := add_mu_information s.(mu_ledger) mu_pdiscover_cost in
            Some {| partition := s.(partition);
                    mu_ledger := mu';
                    pc := S s.(pc);
                    halted := false;
                    result := s.(result);
                    program := s.(program) |}

        | HALT =>
            (* Halt execution *)
            Some {| partition := s.(partition);
                    mu_ledger := s.(mu_ledger);
                    pc := s.(pc);
                    halted := true;
                    result := s.(result);
                    program := s.(program) |}
        end
    end.

(** =========================================================================
    SECTION 4: MULTI-STEP EXECUTION (RUN FUNCTION)
    =========================================================================
    
    Run function: Execute until halt or fuel exhausted.
    Uses fuel parameter to ensure termination of Coq function.
    
    ========================================================================= *)

(** Multi-step execution with fuel *)
Fixpoint run (fuel : nat) (s : State) : State :=
  match fuel with
  | 0%nat => s  (* Out of fuel *)
  | S fuel' =>
      match step s with
      | None => s  (* Already halted *)
      | Some s' =>
          if s'.(halted) then s'  (* Halt reached *)
          else run fuel' s'  (* Continue *)
      end
  end.

(** =========================================================================
    SECTION 5: μ-UPDATE FUNCTION
    =========================================================================
    
    The μ-update function tracks how μ-cost changes across state transitions.
    This is key for verifying μ-monotonicity (A1.4).
    
    ========================================================================= *)

(** Extract μ-total from state *)
Definition mu_of_state (s : State) : Z :=
  s.(mu_ledger).(mu_total).

(** μ-update: Compute μ-cost increase from state transition *)
Definition mu_update (s s' : State) : Z :=
  mu_of_state s' - mu_of_state s.

(** =========================================================================
    SECTION 6: INVARIANTS (PROPERTIES TO BE PROVEN IN A1.4)
    =========================================================================
    
    Core invariants that characterize the Thiele Machine:
    1. μ-monotonicity: μ never decreases
    2. Partition validity: Partitions remain valid
    3. Polynomial time: Execution completes in polynomial time
    
    ========================================================================= *)

(** Invariant 1: μ-Monotonicity *)
Definition mu_monotonic (s s' : State) : Prop :=
  mu_of_state s' >= mu_of_state s.

(** Invariant 2: Partition Validity 
    A partition is valid if:
    - All regions are disjoint
    - All variable IDs are unique
*)
Fixpoint regions_disjoint (regions : list Region) : Prop :=
  match regions with
  | [] => True
  | r :: rest =>
      (forall v, In v r -> ~exists r', In r' rest /\ In v r') /\
      regions_disjoint rest
  end.

Definition partition_valid (p : Partition) : Prop :=
  partition_valid_b p = true.

(** Invariant 3: Polynomial Time Bound
    For a problem of size n, execution completes in O(n³) steps.
    Note: This is a complexity property that depends on the specific program.
    For well-formed programs, halting is guaranteed with sufficient fuel.
*)
Remark polynomial_time_complexity_note :
  (* Well-formed programs halt in polynomial time *)
  (* This is a meta-property about the semantics *)
  forall (n : nat) (s : State) (prog : Program),
    (* With sufficient fuel, well-formed programs halt *)
    (n > 0)%nat -> True.
Proof.
  intros n s prog Hn.
  exact I.
Qed.

(** =========================================================================
    SECTION 7: CORE THEOREMS (A1.4 - PROVEN)
    =========================================================================
    
    These theorems establish the fundamental properties of the Thiele Machine.
    Task A1.4 requires proving these with Qed.
    
    ========================================================================= *)

(** Theorem 1: μ-Monotonicity
    The μ-cost never decreases during execution.
    This is a fundamental conservation law.
*)
Theorem mu_never_decreases :
  forall (s : State) (s' : State),
    step s = Some s' ->
    mu_monotonic s s'.
Proof.
  intros s s' Hstep.
  unfold mu_monotonic, mu_of_state.
  unfold step in Hstep.
  destruct (halted s) eqn:Hhalted.
  - discriminate Hstep.
  - destruct (nth_error (program s) (pc s)) as [instr|] eqn:Hnth.
    + destruct instr; simpl in Hstep.
      * (* PNEW *)
        destruct (existsb (fun r' : Region => region_eqb r r')
                (map snd (modules (partition s)))) eqn:Hdup.
        -- inversion Hstep; subst; clear Hstep. simpl. apply Z.le_ge. apply Z.le_refl.
        -- destruct (existsb (fun r' : Region => negb (disjoint_b r r'))
                 (map snd (modules (partition s)))) eqn:Hov.
           ++ inversion Hstep; subst; clear Hstep. simpl. apply Z.le_ge. apply Z.le_refl.
           ++ set (p' := add_module (partition s) r).
              destruct (partition_valid_b p') eqn:Hpv.
            ** unfold p' in Hpv.
               rewrite Hpv in Hstep.
               inversion Hstep; subst; clear Hstep.
                  simpl.
                  apply add_mu_operational_mu_total_ge.
                  apply mu_pnew_cost_nonneg.
                ** unfold p' in Hpv.
                  rewrite Hpv in Hstep.
                  inversion Hstep; subst; clear Hstep.
                  simpl. apply Z.le_ge. apply Z.le_refl.
      * (* PSPLIT *)
        set (p' := update_partition_split (partition s) m).
        destruct (partition_valid_b p') eqn:Hpv.
          -- unfold p' in Hpv.
             rewrite Hpv in Hstep.
             inversion Hstep; subst; clear Hstep.
            simpl.
            apply add_mu_operational_mu_total_ge.
            apply mu_psplit_cost_nonneg.
        -- unfold p' in Hpv.
          rewrite Hpv in Hstep.
          inversion Hstep; subst; clear Hstep.
          simpl.
          apply add_mu_operational_mu_total_ge.
          apply mu_psplit_cost_nonneg.
      * (* PMERGE *)
        set (p' := update_partition_merge (partition s) m m0).
        destruct (partition_valid_b p') eqn:Hpv.
          -- unfold p' in Hpv.
             rewrite Hpv in Hstep.
             inversion Hstep; subst; clear Hstep.
            simpl.
            apply add_mu_operational_mu_total_ge.
            apply mu_pmerge_cost_nonneg.
         -- unfold p' in Hpv.
           rewrite Hpv in Hstep.
           inversion Hstep; subst; clear Hstep.
           simpl. apply Z.le_ge. apply Z.le_refl.
      * (* LASSERT *)
        destruct (partition_valid_b (partition s)) eqn:Hpv;
          inversion Hstep; subst; clear Hstep.
        -- simpl.
           apply add_mu_operational_mu_total_ge.
           apply mu_lassert_cost_nonneg.
        -- simpl. apply Z.le_ge. apply Z.le_refl.
      * (* LJOIN *)
        inversion Hstep; subst; clear Hstep.
        simpl.
        apply add_mu_operational_mu_total_ge.
        apply mu_lassert_cost_nonneg.
      * (* MDLACC *)
        inversion Hstep; subst; clear Hstep.
        simpl.
        apply add_mu_operational_mu_total_ge.
        apply mu_mdlacc_cost_nonneg.
      * (* PDISCOVER *)
        inversion Hstep; subst; clear Hstep.
        simpl.
        apply add_mu_information_mu_total_ge.
        apply mu_pdiscover_cost_nonneg.
      * (* XFER *)
        inversion Hstep; subst; clear Hstep.
        simpl.
        apply add_mu_operational_mu_total_ge.
        apply mu_emit_cost_nonneg.
      * (* PYEXEC *)
        inversion Hstep; subst; clear Hstep.
        simpl.
        apply add_mu_operational_mu_total_ge.
        apply mu_lassert_cost_nonneg.
      * (* XOR_LOAD *)
        inversion Hstep; subst; clear Hstep.
        simpl.
        apply add_mu_operational_mu_total_ge.
        apply mu_emit_cost_nonneg.
      * (* XOR_ADD *)
        inversion Hstep; subst; clear Hstep.
        simpl.
        apply add_mu_operational_mu_total_ge.
        apply mu_emit_cost_nonneg.
      * (* XOR_SWAP *)
        inversion Hstep; subst; clear Hstep.
        simpl.
        apply add_mu_operational_mu_total_ge.
        apply mu_emit_cost_nonneg.
      * (* XOR_RANK *)
        inversion Hstep; subst; clear Hstep.
        simpl.
        apply add_mu_operational_mu_total_ge.
        apply mu_emit_cost_nonneg.
      * (* EMIT *)
        inversion Hstep; subst; clear Hstep.
        simpl.
        apply add_mu_operational_mu_total_ge.
        apply mu_emit_cost_nonneg.
      * (* ORACLE_HALTS *)
        inversion Hstep; subst; clear Hstep.
        simpl.
        apply add_mu_information_mu_total_ge.
        apply mu_pdiscover_cost_nonneg.
      * (* HALT *)
        inversion Hstep; subst; clear Hstep.
        simpl. apply Z.le_ge. apply Z.le_refl.
    + inversion Hstep; subst; clear Hstep.
      simpl. apply Z.le_ge. apply Z.le_refl.
Qed.

(** Theorem 2: Partition Validity Preservation
    If a partition is valid before a step, it remains valid after.
    
    Note: This is a structural preservation theorem. For PNEW, we assert
    that adding a module maintains validity as a design invariant.
*)
(** Theorem 2: Partition State Preservation
    For computational instructions (non-partition ops), partition structure is preserved.
*)
Theorem partition_preserved_computational :
  forall (s : State) (s' : State) (instr : Instruction),
    nth_error s.(program) s.(pc) = Some instr ->
    s.(halted) = false ->
    step s = Some s' ->
    (forall r, instr <> PNEW r) ->
    (forall m, instr <> PSPLIT m) ->
    (forall m1 m2, instr <> PMERGE m1 m2) ->
    s'.(partition) = s.(partition).
Proof.
  intros s s' instr Hnth Hhalted Hstep Hnot_pnew Hnot_psplit Hnot_pmerge.
  unfold step in Hstep.
  rewrite Hhalted in Hstep.
  rewrite Hnth in Hstep.
  destruct instr.
  - (* PNEW *)
    exfalso. eapply Hnot_pnew. reflexivity.
  - (* PSPLIT *)
    exfalso. eapply Hnot_psplit. reflexivity.
  - (* PMERGE *)
    exfalso. eapply Hnot_pmerge. reflexivity.
  - (* LASSERT *)
    simpl in Hstep. destruct (partition_valid_b (partition s)); injection Hstep as Hstep; subst s'; reflexivity.
  - (* LJOIN *)
    injection Hstep as Hstep; subst s'; reflexivity.
  - (* MDLACC *)
    injection Hstep as Hstep; subst s'; reflexivity.
  - (* PDISCOVER *)
    injection Hstep as Hstep; subst s'; reflexivity.
  - (* XFER *)
    injection Hstep as Hstep; subst s'; reflexivity.
  - (* PYEXEC *)
    injection Hstep as Hstep; subst s'; reflexivity.
  - (* XOR_LOAD *)
    injection Hstep as Hstep; subst s'; reflexivity.
  - (* XOR_ADD *)
    injection Hstep as Hstep; subst s'; reflexivity.
  - (* XOR_SWAP *)
    injection Hstep as Hstep; subst s'; reflexivity.
  - (* XOR_RANK *)
    injection Hstep as Hstep; subst s'; reflexivity.
  - (* EMIT *)
    injection Hstep as Hstep; subst s'; reflexivity.
  - (* ORACLE_HALTS *)
    injection Hstep as Hstep; subst s'; reflexivity.
  - (* HALT *)
    injection Hstep as Hstep; subst s'; reflexivity.
Qed.

(** Theorem 2: Partition Validity Preservation
    If a partition is valid before a step, it remains valid after.

    Note: This relies on the strict PNEW semantics above: new regions must be
    disjoint (duplicates are a no-op; partial overlaps halt).
*)
Theorem partition_validity_preserved :
  forall (s s' : State),
    step s = Some s' ->
    partition_valid (partition s) ->
    partition_valid (partition s').
Proof.
  intros s s' Hstep Hvalid.
  unfold partition_valid in *.
  unfold step in Hstep.
  destruct (halted s) eqn:Hhalted.
  - discriminate Hstep.
  - destruct (nth_error (program s) (pc s)) as [instr|] eqn:Hnth.
    + destruct instr; simpl in Hstep;
      try (injection Hstep as Hstep; subst s'; simpl; exact Hvalid).

    * (* PNEW *)
      destruct (existsb (fun r' : Region => region_eqb r r')
                  (map snd (modules (partition s)))) eqn:Hdup.
      -- (* duplicate: partition unchanged *)
        injection Hstep as Hstep; subst s'.
        simpl. exact Hvalid.
      -- destruct (existsb (fun r' : Region => negb (disjoint_b r r'))
                    (map snd (modules (partition s)))) eqn:Hov.
        ++ (* overlap: partition unchanged *)
          injection Hstep as Hstep; subst s'.
          simpl. exact Hvalid.
        ++ (* disjoint: attempt to add; validity is checked in-step *)
          set (p' := add_module (partition s) r).
          destruct (partition_valid_b p') eqn:Hpv.
            ** unfold p' in Hpv.
               rewrite Hpv in Hstep.
               injection Hstep as Hstep; subst s'.
            simpl. exact Hpv.
            ** unfold p' in Hpv.
               rewrite Hpv in Hstep.
               injection Hstep as Hstep; subst s'.
            simpl. exact Hvalid.

    * (* PSPLIT *)
      set (p' := update_partition_split (partition s) m).
      destruct (partition_valid_b p') eqn:Hpv.
        -- unfold p' in Hpv.
           rewrite Hpv in Hstep.
           injection Hstep as Hstep; subst s'.
        simpl. exact Hpv.
        -- unfold p' in Hpv.
           rewrite Hpv in Hstep.
           injection Hstep as Hstep; subst s'.
        simpl. exact Hvalid.

    * (* PMERGE *)
      set (p' := update_partition_merge (partition s) m m0).
      destruct (partition_valid_b p') eqn:Hpv.
        -- unfold p' in Hpv.
           rewrite Hpv in Hstep.
           injection Hstep as Hstep; subst s'.
        simpl. exact Hpv.
        -- unfold p' in Hpv.
           rewrite Hpv in Hstep.
           injection Hstep as Hstep; subst s'.
        simpl. exact Hvalid.

      * (* LASSERT *)
        rewrite Hvalid in Hstep.
        injection Hstep as Hstep; subst s'.
        simpl. exact Hvalid.

   + (* PC out of bounds: partition unchanged *)
    injection Hstep as Hstep; subst s'.
    simpl. exact Hvalid.
Qed.

(** Theorem 3: Multi-step μ-Monotonicity
    μ-monotonicity holds across multiple steps.
*)
Theorem run_mu_monotonic :
  forall (fuel : nat) (s : State),
    mu_of_state (run fuel s) >= mu_of_state s.
Proof.
  induction fuel as [|fuel' IH]; intros s.
  - (* Base case: fuel = 0 *)
    simpl. lia.
  - (* Inductive case: fuel = S fuel' *)
    simpl.
    destruct (step s) as [s'|] eqn:Hstep.
    + (* Step succeeded *)
      destruct (halted s') eqn:Hhalted'.
      * (* Halted after step *)
        assert (Hmono : mu_of_state s' >= mu_of_state s).
        { apply mu_never_decreases. assumption. }
        lia.
      * (* Not halted, continue running *)
        assert (Hmono : mu_of_state s' >= mu_of_state s).
        { apply mu_never_decreases. assumption. }
        assert (IH' := IH s').
        lia.
    + (* Step failed (already halted) *)
      lia.
Qed.

(** =========================================================================
    SECTION 8: COMPLETENESS PROPERTIES
    =========================================================================
    
    Additional properties showing the machine is well-defined and complete.
    
    ========================================================================= *)

(** Property: Step is deterministic *)
Theorem step_deterministic :
  forall (s : State) (s1 s2 : State),
    step s = Some s1 ->
    step s = Some s2 ->
    s1 = s2.
Proof.
  intros s s1 s2 H1 H2.
  rewrite H1 in H2.
  inversion H2.
  reflexivity.
Qed.

(** Property: Halted states cannot step *)
Theorem halted_cannot_step :
  forall (s : State),
    s.(halted) = true ->
    step s = None.
Proof.
  intros s Hhalted.
  unfold step.
  rewrite Hhalted.
  reflexivity.
Qed.

(** Property: Non-halted states with valid PC can step *)
Theorem valid_pc_can_step :
  forall (s : State),
    s.(halted) = false ->
    (s.(pc) < List.length s.(program))%nat ->
    exists s', step s = Some s'.
Proof.
  intros s Hhalted Hpc.
  unfold step.
  rewrite Hhalted.
  destruct (nth_error (program s) (pc s)) as [instr|] eqn:Hnth.
  - (* Valid instruction *)
    destruct instr.
    + (* PNEW *)
      destruct (existsb (fun r' : Region => region_eqb r r')
                (map snd (modules (partition s)))).
      * eexists; reflexivity.
      * destruct (existsb (fun r' : Region => negb (disjoint_b r r'))
                  (map snd (modules (partition s)))).
        -- eexists; reflexivity.
        -- destruct (partition_valid_b (add_module (partition s) r));
             eexists; reflexivity.
    + (* PSPLIT *)
      destruct (partition_valid_b (update_partition_split (partition s) m));
        eexists; reflexivity.
    + (* PMERGE *)
      destruct (partition_valid_b (update_partition_merge (partition s) m m0));
        eexists; reflexivity.
    + (* LASSERT *)
      destruct (partition_valid_b (partition s));
        eexists; reflexivity.
    + (* LJOIN *) eexists; reflexivity.
    + (* MDLACC *) eexists; reflexivity.
    + (* PDISCOVER *) eexists; reflexivity.
    + (* XFER *) eexists; reflexivity.
    + (* PYEXEC *) eexists; reflexivity.
    + (* XOR_LOAD *) eexists; reflexivity.
    + (* XOR_ADD *) eexists; reflexivity.
    + (* XOR_SWAP *) eexists; reflexivity.
    + (* XOR_RANK *) eexists; reflexivity.
    + (* EMIT *) eexists; reflexivity.
    + (* ORACLE_HALTS *) eexists; reflexivity.
    + (* HALT *) eexists; reflexivity.
  - (* This case is impossible given Hpc *)
    (* nth_error returns None only when pc >= length prog *)
    apply nth_error_None in Hnth.
    lia.
Qed.

(** =========================================================================
    SECTION 9: ALIGNMENT WITH OTHER IMPLEMENTATIONS
    =========================================================================
    
    These properties ensure this Coq semantics aligns with:
    - Python VM (thielecpu/vm.py)
    - Verilog RTL (thielecpu/hardware/thiele_cpu.v)
    
    ========================================================================= *)

(** Property: μ-cost formula matches μ-spec v2.0 *)
Remark mu_costs_align_with_spec :
  mu_pnew_cost = 8 /\
  mu_psplit_cost = 16 /\
  mu_pmerge_cost = 12 /\
  mu_pdiscover_cost = 100 /\
  mu_lassert_cost = 20 /\
  mu_mdlacc_cost = 5 /\
  mu_emit_cost = 1.
Proof.
  unfold mu_pnew_cost, mu_psplit_cost, mu_pmerge_cost,
         mu_pdiscover_cost, mu_lassert_cost, mu_mdlacc_cost,
         mu_emit_cost.
  repeat split; reflexivity.
Qed.

(** =========================================================================
    END OF CORE SEMANTICS
    =========================================================================
    
    SUMMARY:
    ✅ Section 1: State Space S - COMPLETE
    ✅ Section 2: Instruction Set - COMPLETE
    ✅ Section 3: Transition System (step) - COMPLETE
    ✅ Section 4: Multi-step Execution (run) - COMPLETE
    ✅ Section 5: μ-Update Function - COMPLETE
    ✅ Section 6: Invariant Definitions - COMPLETE
    ✅ Section 7: Core Theorems - PARTIALLY COMPLETE
       - μ-Monotonicity: ✅ PROVEN (Qed)
       - Multi-step μ-Monotonicity: ✅ PROVEN (Qed)
       - Partition Validity: ⚠️ ADMITTED (requires more work)
    ✅ Section 8: Completeness Properties - COMPLETE
    ✅ Section 9: Alignment Properties - COMPLETE
    
    NEXT STEPS (A1.4 continuation):
    1. Complete partition_validity_preserved proof
    2. Prove polynomial time bounds (or refine axiom)
    3. Add additional helper lemmas for complex proofs
    
    ========================================================================= *)

(** =========================================================================
    SECTION 10: μ-LEDGER INDEPENDENCE
    =========================================================================
    
    Key property for gauge symmetry: step function's observable behavior
    (partition, pc, halted, result, program) depends only on observable
    components of input state, not on μ-ledger.
    
    ========================================================================= *)

Lemma step_mu_independent : forall s1 s2 s1',
  s1.(partition) = s2.(partition) ->
  s1.(pc) = s2.(pc) ->
  s1.(halted) = s2.(halted) ->
  s1.(result) = s2.(result) ->
  s1.(program) = s2.(program) ->
  step s1 = Some s1' ->
  exists s2',
    step s2 = Some s2' /\
    s1'.(partition) = s2'.(partition) /\
    s1'.(pc) = s2'.(pc) /\
    s1'.(halted) = s2'.(halted) /\
    s1'.(result) = s2'.(result) /\
    s1'.(program) = s2'.(program).
Proof.
  intros s1 s2 s1' Hpart Hpc Hhalt Hres Hprog Hstep1.
  unfold step in *.
  
  (* Rewrite s2 fields to match s1 *)
  unfold step in Hstep1.
  destruct (halted s1) eqn:Hhalt1; [inversion Hstep1 |].
  destruct (nth_error (program s1) (pc s1)) as [i|] eqn:Hinstr1.
  2: { (* nth_error = None → halts *) 
    inversion Hstep1; subst.
    (* Need to show step s2 = Some (halt state) *)
    exists {| partition := partition s2;
              mu_ledger := mu_ledger s2;
              pc := pc s2;
              halted := true;
              result := result s2;
              program := program s2 |}.
    split.
    { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog, Hinstr1. reflexivity. }
    { repeat split; try (rewrite <- Hpart); try (rewrite <- Hpc); try (rewrite <- Hres); try (rewrite <- Hprog); reflexivity. }
  }
  
  (* Case on instruction - construct witness using s1 observables, s2 mu *)
  destruct i as [r | mid | m1 m2 | | | m | | | | | | | | n | | ].
  
  (* PNEW r: branches depend on partition *)
  - (* Case split on the conditions in step s1 *)
    destruct (existsb (fun r' => region_eqb r r') (map snd (modules (partition s1)))) eqn:Hex.
    + (* Exact duplicate: no-op. Return state preserves all observables *)
      (* Construct s2' witness using s1 observable fields (which equal s2's by hypotheses) *)
      exists {| partition := partition s1; mu_ledger := mu_ledger s2; 
                pc := S (pc s1); halted := false; result := result s1; program := program s1 |}.
      split.
      { (* Prove step s2 = Some s2' *)
        unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog, <- Hres. simpl. rewrite Hinstr1. simpl.
        rewrite <- Hpart. simpl. rewrite Hex. simpl. reflexivity.
      }
      { (* Prove observables equal to s1' *)
        injection Hstep1 as Hs1'_eq. subst s1'.
        simpl. split; [reflexivity | split; [reflexivity | split; [reflexivity | 
        split; [reflexivity | reflexivity]]]].
      }
    + (* Exact duplicate false branch - partial overlap check *)
      destruct (existsb (fun r' => negb (disjoint_b r r')) (map snd (modules (partition s1)))) eqn:Hover.
      * (* Partial overlap: halt *)
        exists {| partition := partition s1; mu_ledger := mu_ledger s2; 
                  pc := pc s1; halted := true; result := None; program := program s1 |}.
        split.
        { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog. simpl. rewrite Hinstr1. simpl.
          rewrite <- Hpart. simpl. rewrite Hex, Hover. simpl. reflexivity. }
        { injection Hstep1 as Hs1'_eq. subst s1'.
          simpl. repeat split; reflexivity. }
      * (* No overlap - attempt to add module *)
        destruct (partition_valid_b (add_module (partition s1) r)) eqn:Hvalid.
        -- (* Valid: add module with μ cost *)
           exists {| partition := add_module (partition s1) r; 
                     mu_ledger := add_mu_operational (mu_ledger s2) mu_pnew_cost; 
                     pc := S (pc s1); halted := false; result := result s1; program := program s1 |}.
           split.
           { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog, <- Hres. simpl. rewrite Hinstr1. simpl.
             rewrite <- Hpart. simpl. rewrite Hex, Hover, Hvalid. simpl. reflexivity. }
           { injection Hstep1 as Hs1'_eq. subst s1'.
             simpl. split; [reflexivity | split; [reflexivity | split; [reflexivity | 
             split; [reflexivity | reflexivity]]]]. }
        -- (* Invalid: halt without μ cost *)
           exists {| partition := partition s1; mu_ledger := mu_ledger s2; 
                     pc := pc s1; halted := true; result := None; program := program s1 |}.
           split.
           { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog. simpl. rewrite Hinstr1. simpl.
             rewrite <- Hpart. simpl. rewrite Hex, Hover, Hvalid. simpl. reflexivity. }
           { injection Hstep1 as Hs1'_eq. subst s1'.
             simpl. repeat split; reflexivity. }
  
  (* PSPLIT mid: split module instruction *)
  - destruct (partition_valid_b (update_partition_split (partition s1) mid)) eqn:Hvalid.
    + (* Valid split *)
      exists {| partition := update_partition_split (partition s1) mid;
                mu_ledger := add_mu_operational (mu_ledger s2) mu_psplit_cost;
                pc := S (pc s1); halted := false; result := result s1; program := program s1 |}.
      split.
      { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog, <- Hres. simpl. rewrite Hinstr1. simpl.
        rewrite <- Hpart. simpl. rewrite Hvalid. simpl. reflexivity. }
      { injection Hstep1 as Hs1'_eq. subst s1'.
        simpl. split; [reflexivity | split; [reflexivity | split; [reflexivity | 
        split; [reflexivity | reflexivity]]]]. }
    + (* Invalid split: halt *)
      exists {| partition := partition s1;
                mu_ledger := add_mu_operational (mu_ledger s2) mu_psplit_cost;
                pc := pc s1; halted := true; result := None; program := program s1 |}.
      split.
      { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog. simpl. rewrite Hinstr1. simpl.
        rewrite <- Hpart. simpl. rewrite Hvalid. simpl. reflexivity. }
      { injection Hstep1 as Hs1'_eq. subst s1'.
        simpl. repeat split; reflexivity. }
  
  (* PMERGE m1 m2: merge modules instruction *)
  - destruct (partition_valid_b (update_partition_merge (partition s1) m1 m2)) eqn:Hvalid.
    + (* Valid merge *)
      exists {| partition := update_partition_merge (partition s1) m1 m2;
                mu_ledger := add_mu_operational (mu_ledger s2) mu_pmerge_cost;
                pc := S (pc s1); halted := false; result := result s1; program := program s1 |}.
      split.
      { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog, <- Hres. simpl. rewrite Hinstr1. simpl.
        rewrite <- Hpart. simpl. rewrite Hvalid. simpl. reflexivity. }
      { injection Hstep1 as Hs1'_eq. subst s1'.
        simpl. split; [reflexivity | split; [reflexivity | split; [reflexivity | 
        split; [reflexivity | reflexivity]]]]. }
    + (* Invalid merge: halt *)
      exists {| partition := partition s1; mu_ledger := mu_ledger s2;
                pc := pc s1; halted := true; result := None; program := program s1 |}.
      split.
      { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog. simpl. rewrite Hinstr1. simpl.
        rewrite <- Hpart. simpl. rewrite Hvalid. simpl. reflexivity. }
      { injection Hstep1 as Hs1'_eq. subst s1'.
        simpl. repeat split; reflexivity. }
  
  (* LASSERT: logical assertion instruction *)
  - destruct (partition_valid_b (partition s1)) eqn:Hvalid.
    + (* Assertion passes *)
      exists {| partition := partition s1;
                mu_ledger := add_mu_operational (mu_ledger s2) mu_lassert_cost;
                pc := S (pc s1); halted := false; result := result s1; program := program s1 |}.
      split.
      { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog, <- Hres. simpl. rewrite Hinstr1. simpl.
        rewrite <- Hpart. rewrite Hvalid. simpl. reflexivity. }
      { injection Hstep1 as Hs1'_eq. subst s1'.
        simpl. split; [reflexivity | split; [reflexivity | split; [reflexivity | 
        split; [reflexivity | reflexivity]]]]. }
    + (* Assertion fails: halt *)
      exists {| partition := partition s1; mu_ledger := mu_ledger s2;
                pc := pc s1; halted := true; result := None; program := program s1 |}.
      split.
      { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog. simpl. rewrite Hinstr1. simpl.
        rewrite <- Hpart. rewrite Hvalid. simpl. reflexivity. }
      { injection Hstep1 as Hs1'_eq. subst s1'.
        simpl. repeat split; reflexivity. }
  
  (* LJOIN: logical join instruction *)
  - exists {| partition := partition s1;
              mu_ledger := add_mu_operational (mu_ledger s2) mu_lassert_cost;
              pc := S (pc s1); halted := false; result := result s1; program := program s1 |}.
    split.
    { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog, <- Hres. simpl. rewrite Hinstr1. simpl.
      rewrite <- Hpart. simpl. reflexivity. }
    { injection Hstep1 as Hs1'_eq. subst s1'.
      simpl. split; [reflexivity | split; [reflexivity | split; [reflexivity | 
      split; [reflexivity | reflexivity]]]]. }
  
  (* MDLACC mid: MDL accumulation instruction *)
  - exists {| partition := partition s1;
              mu_ledger := add_mu_operational (mu_ledger s2) mu_mdlacc_cost;
              pc := S (pc s1); halted := false; result := result s1; program := program s1 |}.
    split.
    { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog, <- Hres. simpl. rewrite Hinstr1. simpl.
      rewrite <- Hpart. simpl. reflexivity. }
    { injection Hstep1 as Hs1'_eq. subst s1'.
      simpl. split; [reflexivity | split; [reflexivity | split; [reflexivity | 
      split; [reflexivity | reflexivity]]]]. }
  
  (* PDISCOVER: partition discovery instruction *)
  - exists {| partition := partition s1;
              mu_ledger := add_mu_information (mu_ledger s2) mu_pdiscover_cost;
              pc := S (pc s1); halted := false; result := result s1; program := program s1 |}.
    split.
    { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog, <- Hres. simpl. rewrite Hinstr1. simpl.
      rewrite <- Hpart. simpl. reflexivity. }
    { injection Hstep1 as Hs1'_eq. subst s1'.
      simpl. split; [reflexivity | split; [reflexivity | split; [reflexivity | 
      split; [reflexivity | reflexivity]]]]. }
  
  (* XFER: transfer instruction *)
  - exists {| partition := partition s1;
              mu_ledger := add_mu_operational (mu_ledger s2) mu_emit_cost;
              pc := S (pc s1); halted := false; result := result s1; program := program s1 |}.
    split.
    { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog, <- Hres. simpl. rewrite Hinstr1. simpl.
      rewrite <- Hpart. simpl. reflexivity. }
    { injection Hstep1 as Hs1'_eq. subst s1'.
      simpl. split; [reflexivity | split; [reflexivity | split; [reflexivity | 
      split; [reflexivity | reflexivity]]]]. }
  
  (* PYEXEC: Python execution instruction *)
  - exists {| partition := partition s1;
              mu_ledger := add_mu_operational (mu_ledger s2) mu_lassert_cost;
              pc := S (pc s1); halted := false; result := result s1; program := program s1 |}.
    split.
    { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog, <- Hres. simpl. rewrite Hinstr1. simpl.
      rewrite <- Hpart. simpl. reflexivity. }
    { injection Hstep1 as Hs1'_eq. subst s1'.
      simpl. split; [reflexivity | split; [reflexivity | split; [reflexivity | 
      split; [reflexivity | reflexivity]]]]. }
  
  (* XOR_LOAD: XOR load instruction *)
  - exists {| partition := partition s1;
              mu_ledger := add_mu_operational (mu_ledger s2) mu_emit_cost;
              pc := S (pc s1); halted := false; result := result s1; program := program s1 |}.
    split.
    { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog, <- Hres. simpl. rewrite Hinstr1. simpl.
      rewrite <- Hpart. simpl. reflexivity. }
    { injection Hstep1 as Hs1'_eq. subst s1'.
      simpl. split; [reflexivity | split; [reflexivity | split; [reflexivity | 
      split; [reflexivity | reflexivity]]]]. }
  
  (* XOR_ADD: XOR add instruction *)
  - exists {| partition := partition s1;
              mu_ledger := add_mu_operational (mu_ledger s2) mu_emit_cost;
              pc := S (pc s1); halted := false; result := result s1; program := program s1 |}.
    split.
    { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog, <- Hres. simpl. rewrite Hinstr1. simpl.
      rewrite <- Hpart. simpl. reflexivity. }
    { injection Hstep1 as Hs1'_eq. subst s1'.
      simpl. split; [reflexivity | split; [reflexivity | split; [reflexivity | 
      split; [reflexivity | reflexivity]]]]. }
  
  (* XOR_SWAP: XOR swap instruction *)
  - exists {| partition := partition s1;
              mu_ledger := add_mu_operational (mu_ledger s2) mu_emit_cost;
              pc := S (pc s1); halted := false; result := result s1; program := program s1 |}.
    split.
    { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog, <- Hres. simpl. rewrite Hinstr1. simpl.
      rewrite <- Hpart. simpl. reflexivity. }
    { injection Hstep1 as Hs1'_eq. subst s1'.
      simpl. split; [reflexivity | split; [reflexivity | split; [reflexivity | 
      split; [reflexivity | reflexivity]]]]. }
  
  (* XOR_RANK: XOR rank instruction *)
  - exists {| partition := partition s1;
              mu_ledger := add_mu_operational (mu_ledger s2) mu_emit_cost;
              pc := S (pc s1); halted := false; result := result s1; program := program s1 |}.
    split.
    { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog, <- Hres. simpl. rewrite Hinstr1. simpl.
      rewrite <- Hpart. simpl. reflexivity. }
    { injection Hstep1 as Hs1'_eq. subst s1'.
      simpl. split; [reflexivity | split; [reflexivity | split; [reflexivity | 
      split; [reflexivity | reflexivity]]]]. }
  
  (* EMIT n: emit result instruction *)
  - exists {| partition := partition s1;
              mu_ledger := add_mu_operational (mu_ledger s2) mu_emit_cost;
              pc := S (pc s1); halted := false; result := Some n; program := program s1 |}.
    split.
    { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog. simpl. rewrite Hinstr1. simpl.
      rewrite <- Hpart. simpl. reflexivity. }
    { injection Hstep1 as Hs1'_eq. subst s1'.
      simpl. split; [reflexivity | split; [reflexivity | split; [reflexivity | 
      split; [reflexivity | reflexivity]]]]. }
  
  (* ORACLE_HALTS: oracle halting instruction *)
  - exists {| partition := partition s1;
              mu_ledger := add_mu_information (mu_ledger s2) mu_pdiscover_cost;
              pc := S (pc s1); halted := false; result := result s1; program := program s1 |}.
    split.
    { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog, <- Hres. simpl. rewrite Hinstr1. simpl.
      rewrite <- Hpart. simpl. reflexivity. }
    { injection Hstep1 as Hs1'_eq. subst s1'.
      simpl. split; [reflexivity | split; [reflexivity | split; [reflexivity | 
      split; [reflexivity | reflexivity]]]]. }
  
  (* HALT: halt instruction *)
  - exists {| partition := partition s1; mu_ledger := mu_ledger s2;
              pc := pc s1; halted := true; result := result s1; program := program s1 |}.
    split.
    { unfold step. rewrite <- Hhalt, <- Hpc, <- Hprog, <- Hres. simpl. rewrite Hinstr1. simpl.
      rewrite <- Hpart. simpl. reflexivity. }
    { injection Hstep1 as Hs1'_eq. subst s1'.
      simpl. split; [reflexivity | split; [reflexivity | split; [reflexivity | 
      split; [reflexivity | reflexivity]]]]. }
Qed.

(** Helper lemmas for μ-ledger arithmetic *)
Lemma add_mu_operational_total : forall l delta,
  mu_total (add_mu_operational l delta) = mu_total l + delta.
Proof.
  intros. unfold add_mu_operational. simpl. reflexivity.
Qed.

Lemma add_mu_information_total : forall l delta,
  mu_total (add_mu_information l delta) = mu_total l + delta.
Proof.
  intros. unfold add_mu_information. simpl. reflexivity.
Qed.

(** Corollary: μ-cost deltas are equal for gauge-equivalent states *)
Lemma step_mu_delta_equal : forall s1 s2 s1' s2',
  s1.(partition) = s2.(partition) ->
  s1.(pc) = s2.(pc) ->
  s1.(halted) = s2.(halted) ->
  s1.(result) = s2.(result) ->
  s1.(program) = s2.(program) ->
  step s1 = Some s1' ->
  step s2 = Some s2' ->
  mu_total s1'.(mu_ledger) - mu_total s1.(mu_ledger) =
  mu_total s2'.(mu_ledger) - mu_total s2.(mu_ledger).
Proof.
  intros s1 s2 s1' s2' Hpart Hpc Hhalt Hres Hprog Hstep1 Hstep2.
  (* Use step_mu_independent to relate s1' and a hypothetical s2' from stepping s2 *)
  (* Since s1 and s2 are gauge-equivalent, step_mu_independent gives us that
     the stepped states preserve observable equality. The key is that each
     instruction adds a fixed μ-cost that doesn't depend on initial μ_ledger. *)
  
  (* Unfold step to examine the instruction being executed *)
  unfold step in *.
  destruct (halted s1) eqn:Hhalt1.
  { (* s1 already halted - step returns None, contradicts Hstep1 *)
    try rewrite Hhalt1 in Hstep1; simpl in Hstep1; discriminate. }
  rewrite Hhalt in Hhalt1.
  destruct (halted s2) eqn:Hhalt2.
  { (* s2 already halted - step returns None, contradicts Hstep2 *)
    try rewrite Hhalt2 in Hstep2; simpl in Hstep2; discriminate. }
  
  destruct (nth_error (program s1) (pc s1)) as [i|] eqn:Hinstr1.
  - assert (Hinstr2: nth_error (program s2) (pc s2) = Some i) by (rewrite <- Hprog, <- Hpc, Hinstr1; reflexivity).
    rewrite Hinstr2 in Hstep2.
    (* Now both s1 and s2 execute the same instruction i *)
    (* Each instruction adds a fixed μ-cost, so deltas are equal *)
    destruct i as [r | mid | m1 m2 | | | m | | | | | | | | n | |].
  
    + (* PNEW r *)
    simpl in Hstep1, Hstep2.
    destruct (existsb (fun r' => region_eqb r r') (map snd (modules (partition s1)))) eqn:Hexact1;
    destruct (existsb (fun r' => region_eqb r r') (map snd (modules (partition s2)))) eqn:Hexact2.
    * (* Exact duplicate - no mu change for both *)
      injection Hstep1 as Eq1; injection Hstep2 as Eq2.
      rewrite <- Eq1, <- Eq2; simpl; ring.
    * (* s1 duplicate, s2 not - impossible due to Hpart *)
      exfalso.
      assert (Hexact :
        existsb (fun r' => region_eqb r r') (map snd (modules (partition s1))) =
        existsb (fun r' => region_eqb r r') (map snd (modules (partition s2)))) by (rewrite Hpart; reflexivity).
      rewrite Hexact1 in Hexact; rewrite Hexact2 in Hexact; discriminate.
    * (* s1 not duplicate, s2 is - impossible due to Hpart *)
      exfalso.
      assert (Hexact :
        existsb (fun r' => region_eqb r r') (map snd (modules (partition s1))) =
        existsb (fun r' => region_eqb r r') (map snd (modules (partition s2)))) by (rewrite Hpart; reflexivity).
      rewrite Hexact1 in Hexact; rewrite Hexact2 in Hexact; discriminate.
    * (* Neither is exact duplicate, check partial overlap *)
      destruct (existsb (fun r' => negb (disjoint_b r r')) (map snd (modules (partition s1)))) eqn:Hoverlap1;
      destruct (existsb (fun r' => negb (disjoint_b r r')) (map snd (modules (partition s2)))) eqn:Hoverlap2;
      [ (* Partial overlap - halt, no mu change for both *)
        injection Hstep1 as Eq1; injection Hstep2 as Eq2;
        rewrite <- Eq1, <- Eq2; simpl; ring
      | (* s1 overlaps, s2 doesn't - impossible *)
        exfalso;
        assert (Hoverlap :
          existsb (fun r' => negb (disjoint_b r r')) (map snd (modules (partition s1))) =
          existsb (fun r' => negb (disjoint_b r r')) (map snd (modules (partition s2)))) by (rewrite Hpart; reflexivity);
        rewrite Hoverlap1 in Hoverlap; rewrite Hoverlap2 in Hoverlap; discriminate
      | (* s1 doesn't overlap, s2 does - impossible *)
        exfalso;
        assert (Hoverlap :
          existsb (fun r' => negb (disjoint_b r r')) (map snd (modules (partition s1))) =
          existsb (fun r' => negb (disjoint_b r r')) (map snd (modules (partition s2)))) by (rewrite Hpart; reflexivity);
        rewrite Hoverlap1 in Hoverlap; rewrite Hoverlap2 in Hoverlap; discriminate
      | (* No overlap for either, check partition_valid_b *)
        destruct (partition_valid_b (add_module (partition s1) r)) eqn:Hvalid1;
        destruct (partition_valid_b (add_module (partition s2) r)) eqn:Hvalid2;
        [ (* Valid partition for both - add mu_pnew_cost *)
          injection Hstep1 as Eq1; injection Hstep2 as Eq2;
          rewrite <- Eq1, <- Eq2; simpl mu_ledger;
          rewrite !add_mu_operational_total; ring
        | (* s1 valid, s2 invalid - impossible *)
          assert (Heqvalid: partition_valid_b (add_module (partition s1) r) =
                             partition_valid_b (add_module (partition s2) r)) by (rewrite Hpart; reflexivity);
          rewrite Hvalid1 in Heqvalid; rewrite Hvalid2 in Heqvalid; discriminate
        | (* s1 invalid, s2 valid - impossible *)
          assert (Heqvalid: partition_valid_b (add_module (partition s1) r) =
                             partition_valid_b (add_module (partition s2) r)) by (rewrite Hpart; reflexivity);
          rewrite Hvalid1 in Heqvalid; rewrite Hvalid2 in Heqvalid; discriminate
        | (* Invalid partition for both - halt, no mu change *)
          injection Hstep1 as Eq1; injection Hstep2 as Eq2;
          rewrite <- Eq1, <- Eq2; simpl; ring
        ]
      ].
  
    + (* PSPLIT mid *)
    simpl in Hstep1, Hstep2.
    destruct (partition_valid_b (update_partition_split (partition s1) mid)) eqn:Heqsplit1;
    destruct (partition_valid_b (update_partition_split (partition s2) mid)) eqn:Heqsplit2.
    * (* Valid split for both - add mu_psplit_cost *)
      injection Hstep1 as Eq1; injection Hstep2 as Eq2.
      rewrite <- Eq1, <- Eq2; simpl mu_ledger; rewrite !add_mu_operational_total; ring.
    * (* s1 valid, s2 invalid - impossible *)
      assert (Heqvalid: partition_valid_b (update_partition_split (partition s1) mid) =
                         partition_valid_b (update_partition_split (partition s2) mid)) by (rewrite Hpart; reflexivity).
      rewrite Heqsplit1 in Heqvalid; rewrite Heqsplit2 in Heqvalid; discriminate.
    * (* s1 invalid, s2 valid - impossible *)
      assert (Heqvalid: partition_valid_b (update_partition_split (partition s1) mid) =
                         partition_valid_b (update_partition_split (partition s2) mid)) by (rewrite Hpart; reflexivity).
      rewrite Heqsplit1 in Heqvalid; rewrite Heqsplit2 in Heqvalid; discriminate.
    * (* Invalid split for both - add mu_psplit_cost and halt *)
      injection Hstep1 as Eq1; injection Hstep2 as Eq2.
      rewrite <- Eq1, <- Eq2; simpl mu_ledger; rewrite !add_mu_operational_total; ring.
  
    + (* PMERGE m1 m2 *)
    simpl in Hstep1, Hstep2.
    destruct (partition_valid_b (update_partition_merge (partition s1) m1 m2)) eqn:Heqmerge1;
    destruct (partition_valid_b (update_partition_merge (partition s2) m1 m2)) eqn:Heqmerge2.
    * (* Valid merge for both - add mu_pmerge_cost *)
      injection Hstep1 as Eq1; injection Hstep2 as Eq2.
      rewrite <- Eq1, <- Eq2; simpl mu_ledger; rewrite !add_mu_operational_total; ring.
    * (* s1 valid, s2 invalid - impossible *)
      assert (Heqvalid: partition_valid_b (update_partition_merge (partition s1) m1 m2) =
                         partition_valid_b (update_partition_merge (partition s2) m1 m2)) by (rewrite Hpart; reflexivity).
      rewrite Heqmerge1 in Heqvalid; rewrite Heqmerge2 in Heqvalid; discriminate.
    * (* s1 invalid, s2 valid - impossible *)
      assert (Heqvalid: partition_valid_b (update_partition_merge (partition s1) m1 m2) =
                         partition_valid_b (update_partition_merge (partition s2) m1 m2)) by (rewrite Hpart; reflexivity).
      rewrite Heqmerge1 in Heqvalid; rewrite Heqmerge2 in Heqvalid; discriminate.
    * (* Invalid merge for both - halt, no mu change *)
      injection Hstep1 as Eq1; injection Hstep2 as Eq2.
      rewrite <- Eq1, <- Eq2; simpl; ring.
  
    + (* LASSERT *)
    simpl in Hstep1, Hstep2.
    destruct (partition_valid_b (partition s1)) eqn:Heqassert1;
    destruct (partition_valid_b (partition s2)) eqn:Heqassert2.
    * (* Valid for both *)
      injection Hstep1 as Eq1; injection Hstep2 as Eq2.
      rewrite <- Eq1, <- Eq2; simpl mu_ledger; rewrite !add_mu_operational_total; ring.
    * (* s1 valid, s2 invalid - impossible *)
      assert (Heqvalid: partition_valid_b (partition s1) = partition_valid_b (partition s2)) by (rewrite Hpart; reflexivity).
      rewrite Heqassert1 in Heqvalid; rewrite Heqassert2 in Heqvalid; discriminate.
    * (* s1 invalid, s2 valid - impossible *)
      assert (Heqvalid: partition_valid_b (partition s1) = partition_valid_b (partition s2)) by (rewrite Hpart; reflexivity).
      rewrite Heqassert1 in Heqvalid; rewrite Heqassert2 in Heqvalid; discriminate.
    * (* Invalid for both - halt, no mu change *)
      injection Hstep1 as Eq1; injection Hstep2 as Eq2.
      rewrite <- Eq1, <- Eq2; simpl; ring.
  
    + (* LJOIN *)
    simpl in Hstep1, Hstep2.
    injection Hstep1 as Eq1; injection Hstep2 as Eq2.
    rewrite <- Eq1, <- Eq2; simpl mu_ledger; rewrite !add_mu_operational_total; ring.
  
    + (* MDLACC m *)
    simpl in Hstep1, Hstep2.
    injection Hstep1 as Eq1; injection Hstep2 as Eq2.
    rewrite <- Eq1, <- Eq2; simpl mu_ledger; rewrite !add_mu_operational_total; ring.
  
    + (* PDISCOVER *)
    simpl in Hstep1, Hstep2.
    injection Hstep1 as Eq1; injection Hstep2 as Eq2.
    rewrite <- Eq1, <- Eq2; simpl mu_ledger; rewrite !add_mu_information_total; ring.
  
    + (* XFER *)
    simpl in Hstep1, Hstep2.
    injection Hstep1 as Eq1; injection Hstep2 as Eq2.
    rewrite <- Eq1, <- Eq2; simpl mu_ledger; rewrite !add_mu_operational_total; ring.
  
    + (* PYEXEC *)
    simpl in Hstep1, Hstep2.
    injection Hstep1 as Eq1; injection Hstep2 as Eq2.
    rewrite <- Eq1, <- Eq2; simpl mu_ledger; rewrite !add_mu_operational_total; ring.
  
    + (* XOR_LOAD *)
    simpl in Hstep1, Hstep2.
    injection Hstep1 as Eq1; injection Hstep2 as Eq2.
    rewrite <- Eq1, <- Eq2; simpl mu_ledger; rewrite !add_mu_operational_total; ring.
  
    + (* XOR_ADD *)
    simpl in Hstep1, Hstep2.
    injection Hstep1 as Eq1; injection Hstep2 as Eq2.
    rewrite <- Eq1, <- Eq2; simpl mu_ledger; rewrite !add_mu_operational_total; ring.
  
    + (* XOR_SWAP *)
    simpl in Hstep1, Hstep2.
    injection Hstep1 as Eq1; injection Hstep2 as Eq2.
    rewrite <- Eq1, <- Eq2; simpl mu_ledger; rewrite !add_mu_operational_total; ring.
  
    + (* XOR_RANK *)
    simpl in Hstep1, Hstep2.
    injection Hstep1 as Eq1; injection Hstep2 as Eq2.
    rewrite <- Eq1, <- Eq2; simpl mu_ledger; rewrite !add_mu_operational_total; ring.
  
    + (* EMIT n *)
    simpl in Hstep1, Hstep2.
    injection Hstep1 as Eq1; injection Hstep2 as Eq2.
    rewrite <- Eq1, <- Eq2; simpl mu_ledger; rewrite !add_mu_operational_total; ring.
  
    + (* ORACLE_HALTS *)
    simpl in Hstep1, Hstep2.
    injection Hstep1 as Eq1; injection Hstep2 as Eq2.
    rewrite <- Eq1, <- Eq2; simpl mu_ledger; rewrite !add_mu_information_total; ring.
  
    + (* HALT - no mu change *)
      simpl in Hstep1, Hstep2.
      inversion Hstep1; inversion Hstep2; subst; simpl; ring.
  - assert (Hinstr2: nth_error (program s2) (pc s2) = None) by (rewrite <- Hprog, <- Hpc, Hinstr1; reflexivity).
    simpl in Hstep1; inversion Hstep1; subst s1'.
    rewrite Hinstr2 in Hstep2; simpl in Hstep2; inversion Hstep2; subst s2'.
    simpl; ring.
Qed.

(** =========================================================================
    END OF CORE SEMANTICS
    ========================================================================= *)
