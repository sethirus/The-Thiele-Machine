// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// Copyright 2025 Devon Thiele
//
// See the LICENSE file in the repository root for full terms.
// ============================================================================
// 🚨 CRITICAL SECURITY WARNING 🚨
// ============================================================================
//
// This hardware implements partition-native computation that could be used for:
// - Large-scale cryptanalysis of public-key cryptographic systems
// - Large-scale computational analysis on classical hardware
// - Undermining digital security infrastructure
//
// ETHICAL USE ONLY:
// - This technology is for defensive security research
// - Do not use for offensive cryptanalysis
// - Contact maintainers for security research applications
//
// ============================================================================

`timescale 1ns / 1ps

module thiele_cpu (
    input wire clk,
    input wire rst_n,

    // External interfaces
    output wire [31:0] cert_addr,
    output wire [31:0] status,
    output wire [31:0] error_code,
    output wire [31:0] partition_ops,
    output wire [31:0] mdl_ops,
    output wire [31:0] info_gain,
    output wire [31:0] mu,  // μ-cost accumulator for isomorphism verification

    // Memory interface
    output wire [31:0] mem_addr,
    output wire [31:0] mem_wdata,
    input wire [31:0] mem_rdata,
    output wire mem_we,
    output wire mem_en,

    // Logic engine interface (for Z3 integration)
    output wire logic_req,
    output wire [31:0] logic_addr,
    input wire logic_ack,
    input wire [31:0] logic_data,

    // Python execution interface
    output wire py_req,
    output wire [31:0] py_code_addr,
    input wire py_ack,
    input wire [31:0] py_result,

    // Instruction memory interface
    input wire [31:0] instr_data,
    output wire [31:0] pc
);

// ============================================================================
// PARAMETERS AND CONSTANTS
// ============================================================================

`ifdef YOSYS_LITE
localparam NUM_MODULES = 4;
localparam REGION_SIZE = 16;
`else
localparam NUM_MODULES = 64;
localparam REGION_SIZE = 1024;
`endif
localparam MAX_MU = 32'hFFFFFFFF;

// Instruction opcodes
// Source of truth is the generated header (regenerated by scripts/forge_artifact.sh).
`include "generated_opcodes.vh"

// CSR addresses
localparam [7:0] CSR_CERT_ADDR = 8'h00;
localparam [7:0] CSR_STATUS    = 8'h01;
localparam [7:0] CSR_ERROR     = 8'h02;
localparam [7:0] CSR_PARTITION_OPS = 8'h03;
localparam [7:0] CSR_MDL_OPS   = 8'h04;
localparam [7:0] CSR_INFO_GAIN = 8'h05;

// ============================================================================
// INTERNAL REGISTERS AND WIRES
// ============================================================================

// Program counter
reg [31:0] pc_reg;

// Control and status registers
reg [31:0] csr_cert_addr;
reg [31:0] csr_status;
reg [31:0] csr_error;

// μ-bit accumulator (Q16.16 format)
reg [31:0] mu_accumulator;

// Temporary register for deterministic μ updates in multi-step ops.
reg [31:0] pdiscover_mu_next;

// μ-ALU interface wires
wire [31:0] mu_alu_result;
wire mu_alu_ready;
wire mu_alu_overflow;
reg [2:0] mu_alu_op;
reg [31:0] mu_alu_operand_a;
reg [31:0] mu_alu_operand_b;
reg mu_alu_valid;

// μ-Core interface wires
wire instr_allowed;
wire receipt_required;
wire receipt_accepted;
wire cost_gate_open;
wire partition_gate_open;
wire [31:0] core_status;
wire enforcement_active;
reg [31:0] proposed_cost;
reg [31:0] receipt_value;
reg receipt_valid;

// Temporary registers for task operations
reg [31:0] info_gain_value;

// ---------------------------------------------------------------------------
// Compute state (must mirror Coq-extracted semantics + Python VM)
// ---------------------------------------------------------------------------
reg [31:0] reg_file [0:31];
reg [31:0] data_mem [0:255];

// Performance counters
reg [31:0] partition_ops_counter;
reg [31:0] mdl_ops_counter;
reg [31:0] info_gain_counter;

// Current instruction
wire [31:0] current_instr;
wire [7:0] opcode;
wire [7:0] operand_a;
wire [7:0] operand_b;
wire [7:0] operand_cost;

// Module management
reg [31:0] module_table [0:NUM_MODULES-1];
reg [31:0] region_table [0:NUM_MODULES-1][0:REGION_SIZE-1];
reg [5:0] current_module;
reg [5:0] next_module_id;
reg [31:0] swap_temp;
reg [31:0] rank_temp;

// State machine
reg [3:0] state;
reg [3:0] alu_return_state;  // State to return to after ALU operation
reg [7:0] alu_context;       // Context for ALU operation (which task/phase)

// Loop variables for initialization
reg [31:0] i, j, region_size, even_count, odd_count, size_a, size_b, total_size, module_size, mdl_cost, temp_size, src_size, dest_size;
localparam [3:0] STATE_FETCH = 4'h0;
localparam [3:0] STATE_DECODE = 4'h1;
localparam [3:0] STATE_EXECUTE = 4'h2;
localparam [3:0] STATE_MEMORY = 4'h3;
localparam [3:0] STATE_LOGIC = 4'h4;
localparam [3:0] STATE_PYTHON = 4'h5;
localparam [3:0] STATE_COMPLETE = 4'h6;
localparam [3:0] STATE_ALU_WAIT = 4'h7;        // Wait for μ-ALU operation
localparam [3:0] STATE_ALU_WAIT2 = 4'h8;       // Second ALU wait (for pdiscover)
localparam [3:0] STATE_RECEIPT_HOLD = 4'h9;    // Hold receipt valid for one cycle
localparam [3:0] STATE_PDISCOVER_LAUNCH2 = 4'hA;   // Launch second μ-ALU op for PDISCOVER
localparam [3:0] STATE_PDISCOVER_ARM2 = 4'hB;      // Extra arm cycle before WAIT2 samples μ-ALU

// Context values for ALU operations
localparam [7:0] ALU_CTX_MDLACC = 8'h01;
localparam [7:0] ALU_CTX_PDISCOVER1 = 8'h02;   // First ALU op in pdiscover
localparam [7:0] ALU_CTX_PDISCOVER2 = 8'h03;   // Second ALU op in pdiscover
localparam [7:0] ALU_CTX_ORACLE = 8'h04;

// ============================================================================
// ASSIGNMENTS
// ============================================================================

assign pc = pc_reg;
assign current_instr = instr_data;
assign opcode = current_instr[31:24];
assign operand_a = current_instr[23:16];
assign operand_b = current_instr[15:8];
assign operand_cost = current_instr[7:0];

assign cert_addr = csr_cert_addr;
assign status = csr_status;
assign error_code = csr_error;
assign partition_ops = partition_ops_counter;
assign mdl_ops = mdl_ops_counter;
assign info_gain = info_gain_counter;
assign mu = mu_accumulator;  // Export μ-cost for 3-way isomorphism verification

// ============================================================================
// MAIN CPU LOGIC
// ============================================================================

always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        // Reset logic
        pc_reg <= 32'h0;
        csr_cert_addr <= 32'h0;
        csr_status <= 32'h0;
        csr_error <= 32'h0;
        mu_accumulator <= 32'h0;
        partition_ops_counter <= 32'h0;
        mdl_ops_counter <= 32'h0;
        info_gain_counter <= 32'h0;
        current_module <= 6'h0;
        next_module_id <= 6'h1;
        state <= STATE_FETCH;

`ifndef SYNTHESIS
        // Initialize module table (simulation-only; most synthesis flows cannot
        // implement full memory clears on reset, and Yosys will reject async
        // reset writes to inferred memories).
        for (i = 0; i < NUM_MODULES; i = i + 1) begin
            module_table[i] <= 32'h0;
            for (j = 0; j < REGION_SIZE; j = j + 1) begin
                region_table[i][j] <= 32'h0;
            end
        end

        // Initialize compute state (simulation-only)
        for (i = 0; i < 32; i = i + 1) begin
            reg_file[i] <= 32'h0;
        end
        for (i = 0; i < 256; i = i + 1) begin
            data_mem[i] <= 32'h0;
        end
`endif

    end else begin
        case (state)
            STATE_FETCH: begin
                // Fetch next instruction
                state <= STATE_DECODE;
            end

            STATE_DECODE: begin
                // Decode instruction and calculate proposed μ-cost for μ-Core
                proposed_cost <= mu_accumulator + operand_cost;
                state <= STATE_EXECUTE;
            end

            STATE_EXECUTE: begin
                case (opcode)
                    OPCODE_PNEW: begin
                        // Create new partition module
                        // μ-Core enforcement: check partition gate is open
                        if (instr_allowed && partition_gate_open) begin
                            execute_pnew(operand_a, operand_b);
                            // Coq semantics: vm_mu := s.vm_mu + instruction_cost
                            mu_accumulator <= mu_accumulator + {24'h0, operand_cost};
                            pc_reg <= pc_reg + 4;
                            state <= STATE_FETCH;
                        end else begin
                            // μ-Core denied operation - signal error
                            csr_error <= 32'hA; // MU_CORE_DENIED
                            pc_reg <= pc_reg + 4;
                            state <= STATE_FETCH;
                        end
                    end

                    OPCODE_PSPLIT: begin
                        // Split existing module
                        // μ-Core enforcement: check partition gate is open
                        if (instr_allowed && partition_gate_open) begin
                            execute_psplit(operand_a, operand_b);
                            // Coq semantics: vm_mu := s.vm_mu + instruction_cost
                            mu_accumulator <= mu_accumulator + {24'h0, operand_cost};
                            pc_reg <= pc_reg + 4;
                            state <= STATE_FETCH;
                        end else begin
                            // μ-Core denied operation - signal error
                            csr_error <= 32'hA; // MU_CORE_DENIED
                            pc_reg <= pc_reg + 4;
                            state <= STATE_FETCH;
                        end
                    end

                    OPCODE_PMERGE: begin
                        // Merge two modules
                        // μ-Core enforcement: check partition gate is open
                        if (instr_allowed && partition_gate_open) begin
                            execute_pmerge(operand_a, operand_b);
                            // Coq semantics: vm_mu := s.vm_mu + instruction_cost
                            mu_accumulator <= mu_accumulator + {24'h0, operand_cost};
                            pc_reg <= pc_reg + 4;
                            state <= STATE_FETCH;
                        end else begin
                            // μ-Core denied operation - signal error
                            csr_error <= 32'hA; // MU_CORE_DENIED
                            pc_reg <= pc_reg + 4;
                            state <= STATE_FETCH;
                        end
                    end

                    OPCODE_LASSERT: begin
                        // Logic assertion with proof certificate
                        // Coq semantics: vm_mu := s.vm_mu + instruction_cost
                        //
                        // QUANTITATIVE NO FREE INSIGHT (StateSpaceCounting.v):
                        // operand_cost ≥ String.length(formula) enforced by assembler
                        // This ensures Δμ ≥ formula_bit_length as proven in Coq
                        mu_accumulator <= mu_accumulator + {24'h0, operand_cost};
                        state <= STATE_LOGIC;
                    end

                    OPCODE_LJOIN: begin
                        // Join certificates
                        execute_ljoin(operand_a, operand_b);
                        // Coq semantics: vm_mu := s.vm_mu + instruction_cost
                        mu_accumulator <= mu_accumulator + {24'h0, operand_cost};
                        pc_reg <= pc_reg + 4;
                        state <= STATE_FETCH;
                    end

                    OPCODE_EMIT: begin
                        // Emit value
                        execute_emit(operand_a, operand_b);
                        // Coq semantics: vm_mu := s.vm_mu + instruction_cost
                        mu_accumulator <= mu_accumulator + {24'h0, operand_cost};
                        pc_reg <= pc_reg + 4;
                        state <= STATE_FETCH;
                    end

                    OPCODE_REVEAL: begin
                        // Reveal hidden information (increases mu by specified bits)
                        // This instruction charges μ-cost for revealing previously hidden structural info
                        // 
                        // μ-cost calculation:
                        //   total_cost = instruction_cost + revelation_cost
                        //   instruction_cost = operand_cost (from instruction encoding)
                        //   revelation_cost = operand_a << 8 (Q16.16 fixed point: operand_a * 256)
                        //
                        // operand_a: number of bits being revealed (integer)
                        // operand_b: certificate reference (stored in cert_addr CSR)
                        //
                        // Example: Revealing 5 bits costs 5.0 μ-bits in Q16.16 = 5 << 16 = 0x50000
                        //          But operand_a holds 5, so we shift: {16'h0, 5, 8'h0} = 0x00050000
                        //
                        // Coq semantics: vm_mu := s.vm_mu + instruction_cost + (bits * mu_bit_scale)
                        mu_accumulator <= mu_accumulator + {24'h0, operand_cost} + {16'h0, operand_a, 8'h0};
                        csr_cert_addr <= {24'h0, operand_b}; // Store cert reference
                        pc_reg <= pc_reg + 4;
                        state <= STATE_FETCH;
                    end

                    OPCODE_XFER: begin
                        // Transfer data
                        execute_xfer(operand_a, operand_b);
                        // Coq semantics: vm_mu := s.vm_mu + instruction_cost
                        mu_accumulator <= mu_accumulator + {24'h0, operand_cost};
                        pc_reg <= pc_reg + 4;
                        state <= STATE_FETCH;
                    end

                    OPCODE_PYEXEC: begin
                        // Execute Python code
                        // Coq semantics: vm_mu := s.vm_mu + instruction_cost
                        mu_accumulator <= mu_accumulator + {24'h0, operand_cost};
                        state <= STATE_PYTHON;
                    end

                    OPCODE_CHSH_TRIAL: begin
                        // CHSH trial event.
                        // Encoding convention used by the 3-layer CHSH gate:
                        //   operand_a[1:0] = {x,y}
                        //   operand_b[1:0] = {a,b}
                        // Cost byte is reserved for μ-cost and should be 0.
                        // Invalid bit encodings latch an error.
                        if ((operand_a[7:2] != 6'b0) || (operand_b[7:2] != 6'b0)) begin
                            csr_error <= 32'h1;
                        end
                        // Coq semantics: vm_mu := s.vm_mu + instruction_cost
                        mu_accumulator <= mu_accumulator + {24'h0, operand_cost};
                        pc_reg <= pc_reg + 4;
                        state <= STATE_FETCH;
                    end

                    OPCODE_MDLACC: begin
                        // Accumulate MDL for module; operand_a==0 means current module
                        // Note: execute_mdlacc handles state transition to ALU_WAIT
                        if (operand_a == 8'h00) begin
                            execute_mdlacc(current_module);
                        end else begin
                            execute_mdlacc(operand_a);
                        end
                        // Don't set pc_reg or state here - task handles it
                    end

                    OPCODE_PDISCOVER: begin
                        // Partition discovery: compute information gain
                        // Note: execute_pdiscover handles state transition to ALU_WAIT
                        execute_pdiscover(operand_a, operand_b);
                        // Don't set pc_reg or state here - task handles it
                    end

                    OPCODE_XOR_LOAD: begin
                        // Load XOR matrix row
                        execute_xor_load(operand_a, operand_b);
                        // Coq semantics: vm_mu := s.vm_mu + instruction_cost
                        mu_accumulator <= mu_accumulator + {24'h0, operand_cost};
                        pc_reg <= pc_reg + 4;
                        state <= STATE_FETCH;
                    end

                    OPCODE_XOR_ADD: begin
                        // Add rows in XOR matrix
                        execute_xor_add(operand_a, operand_b);
                        // Coq semantics: vm_mu := s.vm_mu + instruction_cost
                        mu_accumulator <= mu_accumulator + {24'h0, operand_cost};
                        pc_reg <= pc_reg + 4;
                        state <= STATE_FETCH;
                    end

                    OPCODE_XOR_SWAP: begin
                        // Swap rows in XOR matrix
                        execute_xor_swap(operand_a, operand_b);
                        // Coq semantics: vm_mu := s.vm_mu + instruction_cost
                        mu_accumulator <= mu_accumulator + {24'h0, operand_cost};
                        pc_reg <= pc_reg + 4;
                        state <= STATE_FETCH;
                    end

                    OPCODE_XOR_RANK: begin
                        // Compute rank of XOR matrix
                        execute_xor_rank(operand_a, operand_b);
                        // Coq semantics: vm_mu := s.vm_mu + instruction_cost
                        mu_accumulator <= mu_accumulator + {24'h0, operand_cost};
                        pc_reg <= pc_reg + 4;
                        state <= STATE_FETCH;
                    end

                    OPCODE_ORACLE_HALTS: begin
                        // Hyper-Thiele Oracle Primitive
                        // In hardware, this would trigger an external oracle interface
                        // For now, we simulate the cost and interface
                        // Note: execute_oracle_halts handles state transition to ALU_WAIT
                        execute_oracle_halts(operand_a, operand_b);
                        // Don't set pc_reg or state here - task handles it
                    end

                    OPCODE_HALT: begin
                        // Note: RTL formerly auto-charged MDL here, but this contaminates mu_accumulator
                        // with ALU results. For 3-way isomorphism, HALT must be pure.
                        // If MDL charging is needed, use explicit MDLACC before HALT.
                        // Coq semantics: vm_mu := s.vm_mu + instruction_cost
                        mu_accumulator <= mu_accumulator + {24'h0, operand_cost};
                        pc_reg <= pc_reg + 4;
                        state <= STATE_FETCH;
                    end

                    default: begin
                        // Unknown opcode
                        csr_error <= 32'h1;
                        pc_reg <= pc_reg + 4;
                        state <= STATE_FETCH;
                    end
                endcase
            end

            STATE_LOGIC: begin
                // Handle logic engine operations
                if (logic_ack) begin
                    // Logic operation complete
                    csr_cert_addr <= logic_data;
                    pc_reg <= pc_reg + 4;
                    state <= STATE_FETCH;
                end
            end

            STATE_PYTHON: begin
                // Handle Python execution
                if (py_ack) begin
                    // Python execution complete
                    csr_status <= py_result;
                    pc_reg <= pc_reg + 4;
                    state <= STATE_FETCH;
                end
            end

            STATE_ALU_WAIT: begin
                // Wait for μ-ALU operation to complete
                if (mu_alu_ready) begin
                    mu_alu_valid <= 1'b0;

                    // Handle result based on context
                    case (alu_context)
                        ALU_CTX_MDLACC: begin
                            if (mu_alu_overflow) begin
                                csr_error <= 32'h6; // μ-bit overflow
                                pc_reg <= pc_reg + 4;
                                state <= STATE_FETCH;
                            end else begin
                                $display("MDLACC size=%0d mdl_cost=%0d mu_acc(before)=%0d mu_acc(after)=%0d",
                                        module_size, mdl_cost >> 16, mu_accumulator >> 16, mu_alu_result >> 16);
                                mu_accumulator <= mu_alu_result;
                                csr_status <= 32'h5; // MDL accumulation successful
                                mdl_ops_counter <= mdl_ops_counter + 1;

                                // Provide receipt to μ-Core and transition to hold state
                                receipt_value <= mu_alu_result;
                                receipt_valid <= 1'b1;
                                state <= STATE_RECEIPT_HOLD;
                            end
                        end

                        ALU_CTX_PDISCOVER1: begin
                            if (mu_alu_overflow) begin
                                csr_error <= 32'h8; // Information gain overflow
                                pc_reg <= pc_reg + 4;
                                state <= STATE_FETCH;
                            end else begin
                                info_gain_value <= mu_alu_result;

                                // Accumulate info gain directly. The μ-ALU result is already
                                // in Q16.16; a second μ-ALU transaction here is fragile under
                                // registered ready/result timing and can consume stale values.
                                pdiscover_mu_next = mu_accumulator + mu_alu_result;
                                $display("PDISCOVER info_gain=%0d mu_acc(before)=%0d mu_acc(after)=%0d",
                                        mu_alu_result >> 16, mu_accumulator >> 16, pdiscover_mu_next >> 16);
                                mu_accumulator <= pdiscover_mu_next;
                                csr_status <= 32'h6; // Discovery successful
                                partition_ops_counter <= partition_ops_counter + 1;

                                // Provide receipt to μ-Core and transition to hold state
                                receipt_value <= pdiscover_mu_next;
                                receipt_valid <= 1'b1;
                                state <= STATE_RECEIPT_HOLD;
                            end
                        end

                        ALU_CTX_ORACLE: begin
                            if (mu_alu_overflow) begin
                                csr_error <= 32'h6; // μ-bit overflow
                            end else begin
                                mu_accumulator <= mu_alu_result;
                                csr_status <= 32'h42; // "Answer to Life, Universe, and Everything" placeholder
                                $display("ORACLE_HALTS invoked - Hyper-Thiele transition");
                            end
                            pc_reg <= pc_reg + 4;
                            state <= STATE_FETCH;
                        end

                        default: begin
                            pc_reg <= pc_reg + 4;
                            state <= alu_return_state;
                        end
                    endcase
                end
            end

            STATE_PDISCOVER_LAUNCH2: begin
                // Second-stage PDISCOVER: accumulate the previously computed info gain.
                mu_alu_op <= 3'd0;  // ADD
                mu_alu_operand_a <= mu_accumulator;
                mu_alu_operand_b <= info_gain_value;
                mu_alu_valid <= 1'b1;
                alu_context <= ALU_CTX_PDISCOVER2;
                // Give μ-ALU enough cycles that WAIT2 doesn't consume the
                // previous operation's registered outputs.
                state <= STATE_PDISCOVER_ARM2;
            end

            STATE_PDISCOVER_ARM2: begin
                state <= STATE_ALU_WAIT2;
            end

            STATE_ALU_WAIT2: begin
                // Second ALU wait (for pdiscover)
                if (mu_alu_ready) begin
                    mu_alu_valid <= 1'b0;

                    if (alu_context == ALU_CTX_PDISCOVER2) begin
                        if (mu_alu_overflow) begin
                            csr_error <= 32'h6; // μ-bit overflow
                            pc_reg <= pc_reg + 4;
                            state <= STATE_FETCH;
                        end else begin
                            $display("PDISCOVER info_gain=%0d mu_acc(before)=%0d mu_acc(after)=%0d",
                                    info_gain_value >> 16, mu_accumulator >> 16, mu_alu_result >> 16);
                            mu_accumulator <= mu_alu_result;
                            csr_status <= 32'h6; // Discovery successful
                            partition_ops_counter <= partition_ops_counter + 1;

                            // Provide receipt to μ-Core and transition to hold state
                            receipt_value <= mu_alu_result;
                            receipt_valid <= 1'b1;
                            state <= STATE_RECEIPT_HOLD;
                        end
                    end else begin
                        pc_reg <= pc_reg + 4;
                        state <= alu_return_state;
                    end
                end
            end

            STATE_RECEIPT_HOLD: begin
                // Hold receipt valid for one cycle, then clear
                receipt_valid <= 1'b0;
                pc_reg <= pc_reg + 4;
                state <= STATE_FETCH;
            end

            default: begin
                state <= STATE_FETCH;
            end
        endcase
    end
end

// ============================================================================
// PARTITION OPERATIONS
// ============================================================================

task execute_pnew;
    input [7:0] region_spec_a;
    input [7:0] region_spec_b;
    begin
        // μ-Core enforcement is now checked in STATE_EXECUTE before calling this task.
        // Canonical PNEW encoding used by Python ISA: create/dedup singleton region {operand_a}.
            // operand_b is currently unused (reserved).
            integer found;
            integer found_id;
            found = 0;
            found_id = 0;

            for (i = 0; i < NUM_MODULES; i = i + 1) begin
                if (i < next_module_id) begin
                    if (module_table[i] == 32'd1 && region_table[i][0] == region_spec_a) begin
                        found = 1;
                        found_id = i;
                    end
                end
            end

            if (found) begin
                current_module <= found_id[5:0];
                csr_status <= 32'h1; // Success (dedup)
                $display("PNEW dedup: region={%0d} -> module %0d", region_spec_a, found_id);
            end else if (next_module_id < NUM_MODULES) begin
                module_table[next_module_id] <= 32'd1;
                region_table[next_module_id][0] <= region_spec_a;
                for (i = 1; i < REGION_SIZE; i = i + 1) begin
                    region_table[next_module_id][i] <= 32'h0;
                end
                current_module <= next_module_id;
                next_module_id <= next_module_id + 1;

                csr_status <= 32'h1; // Success
                partition_ops_counter <= partition_ops_counter + 1;
                $display("PNEW new: region={%0d} -> module %0d", region_spec_a, next_module_id);
            end else begin
                csr_error <= 32'h2; // No available modules
            end
    end
endtask

task execute_psplit;
    input [7:0] module_id;
    input [7:0] predicate;
    reg [1:0] pred_mode;
    reg [5:0] pred_param;
    reg [31:0] element_value;
    reg matches_predicate;
    begin
        // Split module based on predicate encoding
        // Predicate format (8 bits):
        //   [7:6] = Mode: 00=even/odd, 01=threshold, 10=bitwise, 11=modulo
        //   [5:0] = Parameter (threshold value, bitmask, or modulo divisor)
        if (module_id < next_module_id && next_module_id < NUM_MODULES - 1) begin
            region_size = module_table[module_id];
            
            pred_mode = predicate[7:6];
            pred_param = predicate[5:0];

            even_count = 0;
            odd_count = 0;

            for (i = 0; i < REGION_SIZE; i = i + 1) begin
                if (i < region_size) begin
                    element_value = region_table[module_id][i];
                    
                    // Evaluate predicate based on mode
                    case (pred_mode)
                        // 00=even/odd: pred_param[0]=0 => even, pred_param[0]=1 => odd
                        2'b00: matches_predicate = (element_value[0] == pred_param[0]);
                        2'b01: matches_predicate = element_value >= pred_param; // Threshold
                        2'b10: matches_predicate = (element_value & (1 << pred_param)) != 0; // Bitwise test
                        // 11=modulo divisibility (synth-safe subset): only supports power-of-two divisors.
                        // divisor = pred_param + 1; if divisor is power-of-two, then (x % divisor)==0 iff (x & (divisor-1))==0.
                        // Here (divisor-1) == pred_param.
                        2'b11: matches_predicate = (((pred_param + 1) & pred_param) == 0) ? ((element_value & pred_param) == 0) : 1'b0;
                        default: matches_predicate = 0;
                    endcase
                    
                    if (matches_predicate) begin
                        region_table[next_module_id][even_count] <= element_value;
                        even_count = even_count + 1;
                    end else begin
                        region_table[next_module_id + 1][odd_count] <= element_value;
                        odd_count = odd_count + 1;
                    end
                end
            end

            module_table[next_module_id] <= even_count;
            module_table[next_module_id + 1] <= odd_count;

            // Coq semantics: graph_psplit replaces module_id with the two new
            // modules; the parent must be removed (no "zombie parent").
            module_table[module_id] <= 32'h0;

            next_module_id <= next_module_id + 2;

            csr_status <= 32'h2; // Split successful
            partition_ops_counter <= partition_ops_counter + 1;
        end else begin
            csr_error <= 32'h3; // Invalid module or no space
        end
    end
endtask

task execute_pmerge;
    input [7:0] module_a;
    input [7:0] module_b;
    begin
        // Merge two modules
        if (module_a < next_module_id && module_b < next_module_id && module_a != module_b) begin
            size_a = module_table[module_a];
            size_b = module_table[module_b];
            total_size = size_a + size_b;

            if (total_size <= REGION_SIZE) begin
                // Copy regions
                for (i = 0; i < REGION_SIZE; i = i + 1) begin
                    if (i < size_a) begin
                        region_table[next_module_id][i] <= region_table[module_a][i];
                    end
                end
                for (i = 0; i < REGION_SIZE; i = i + 1) begin
                    if (i < size_b) begin
                        region_table[next_module_id][i + size_a] <= region_table[module_b][i];
                    end
                end

                module_table[next_module_id] <= total_size;
                module_table[module_a] <= 32'h0; // Mark as free
                module_table[module_b] <= 32'h0; // Mark as free
                current_module <= next_module_id;
                next_module_id <= next_module_id + 1;

                csr_status <= 32'h3; // Merge successful
                partition_ops_counter <= partition_ops_counter + 1;
            end else begin
                csr_error <= 32'h4; // Region too large
            end
        end else begin
            csr_error <= 32'h5; // Invalid modules
        end
    end
endtask

// ============================================================================
// LOGIC AND PYTHON OPERATIONS
// ============================================================================

task execute_ljoin;
    input [7:0] cert_a;
    input [7:0] cert_b;
    begin
        // Join two certificates
        // This would interface with the logic engine
        csr_cert_addr <= {cert_a, cert_b, 16'h0};
        csr_status <= 32'h4; // Join operation
    end
endtask

task execute_mdlacc;
    input [7:0] module_id;
    begin
        // Accumulate μ-bits for MDL cost using Q16.16 arithmetic
        if (module_id < next_module_id) begin
            module_size = module_table[module_id];

            // MDL calculation: partition_bits = bit_length(max_element) * module_size
            if (module_size > 0) begin
                integer max_element;
                integer bit_length;
                integer k;
                max_element = 0;
                // Use constant loop bound for synthesis
                for (k = 0; k < REGION_SIZE; k = k + 1) begin
                    if (k < module_size && region_table[module_id][k] > max_element) begin
                        max_element = region_table[module_id][k];
                    end
                end
                // Compute ceil(log2(max_element + 1)) deterministically.
                // NOTE: Do not depend on combinational clz8_out in the same
                // procedural block after assigning clz8_in; that introduces
                // delta-cycle ordering issues and can produce 'x' in simulation.
                bit_length = ceil_log2_8(max_element + 1);
                // Convert to Q16.16: mdl_cost = (bit_length * module_size) << 16
                mdl_cost = (bit_length * module_size) << 16;
            end else begin
                mdl_cost = 0;
            end

            // Use μ-ALU for Q16.16 addition with saturation
            mu_alu_op <= 3'd0;  // ADD
            mu_alu_operand_a <= mu_accumulator;
            mu_alu_operand_b <= mdl_cost;
            mu_alu_valid <= 1'b1;

            // Set up context and transition to wait state
            alu_context <= ALU_CTX_MDLACC;
            alu_return_state <= STATE_FETCH;
            state <= STATE_ALU_WAIT;
        end else begin
            csr_error <= 32'h7; // Invalid module
        end
    end
endtask

task execute_pdiscover;
    input [7:0] before_count;
    input [7:0] after_count;
    begin
        // Compute information gain: log2(before/after) for partition discovery
        if (before_count > 0 && after_count > 0 && after_count <= before_count) begin
            // Use μ-ALU to compute information gain
            mu_alu_op <= 3'd5;  // INFO_GAIN
            mu_alu_operand_a <= before_count;  // before (integer)
            mu_alu_operand_b <= after_count;   // after (integer)
            mu_alu_valid <= 1'b1;

            // Set up context for first ALU operation
            alu_context <= ALU_CTX_PDISCOVER1;
            alu_return_state <= STATE_FETCH;
            state <= STATE_ALU_WAIT;
        end else begin
            csr_error <= 32'h9; // Invalid discovery parameters
        end
    end
endtask

task execute_emit;
    input [7:0] value_a;
    input [7:0] value_b;
    begin
        // Emit value to output
        // Match Python VM semantics: accumulate value_b into info_gain_counter
        info_gain_counter <= info_gain_counter + value_b;
        csr_status <= {value_a, value_b, 16'h0};
    end
endtask

task execute_xfer;
    input [7:0] dest;
    input [7:0] src;
    begin
        // Register transfer (matches Python VM + Coq kernel semantics)
        reg_file[dest[4:0]] <= reg_file[src[4:0]];
        csr_status <= 32'h6; // Transfer successful
    end
endtask

// ============================================================================
// XOR OPERATIONS
// ============================================================================

task execute_xor_load;
    input [7:0] dest;
    input [7:0] addr;
    begin
        reg_file[dest[4:0]] <= data_mem[addr];
        csr_status <= 32'h7; // XOR load successful
    end
endtask

task execute_xor_add;
    input [7:0] dest;
    input [7:0] src;
    begin
        reg_file[dest[4:0]] <= reg_file[dest[4:0]] ^ reg_file[src[4:0]];
        csr_status <= 32'h8; // XOR add successful
    end
endtask

task execute_xor_swap;
    input [7:0] a;
    input [7:0] b;
    begin
        reg_file[a[4:0]] <= reg_file[b[4:0]];
        reg_file[b[4:0]] <= reg_file[a[4:0]];
        csr_status <= 32'h9; // XOR swap successful
    end
endtask

task execute_xor_rank;
    input [7:0] dest;
    input [7:0] src;
    integer k;
    reg [31:0] v;
    reg [31:0] cnt;
    begin
        v = reg_file[src[4:0]];
        cnt = 0;
        for (k = 0; k < 32; k = k + 1) begin
            cnt = cnt + v[k];
        end
        reg_file[dest[4:0]] <= cnt;
        csr_status <= cnt;
    end
endtask

task execute_oracle_halts;
    input [7:0] desc_ptr_a;
    input [7:0] desc_ptr_b;
    begin
        // Hyper-Thiele Oracle Operation
        // This is a semantic primitive that is not Turing-computable.
        // In a physical realization, this would interface with a hyper-computer
        // or be a placeholder for a non-computable transition.

        // Charge the distinct "Oracle μ" cost (arbitrary high value)
        // Using μ-ALU to add cost
        mu_alu_op <= 3'd0;  // ADD
        mu_alu_operand_a <= mu_accumulator;
        mu_alu_operand_b <= 32'd1000000; // High cost
        mu_alu_valid <= 1'b1;

        // Set up context and transition to wait state
        alu_context <= ALU_CTX_ORACLE;
        alu_return_state <= STATE_FETCH;
        state <= STATE_ALU_WAIT;
    end
endtask

// ============================================================================
// EXTERNAL INTERFACE LOGIC
// ============================================================================

// Instantiate μ-ALU
mu_alu mu_alu_inst (
    .clk(clk),
    .rst_n(rst_n),
    .op(mu_alu_op),
    .operand_a(mu_alu_operand_a),
    .operand_b(mu_alu_operand_b),
    .valid(mu_alu_valid),
    .result(mu_alu_result),
    .ready(mu_alu_ready),
    .overflow(mu_alu_overflow)
);

// Instantiate μ-Core (Partition Isomorphism Enforcement)
mu_core mu_core_inst (
    .clk(clk),
    .rst_n(rst_n),
    .instruction(current_instr),
    .instr_valid(state == STATE_DECODE || state == STATE_EXECUTE),
    .instr_allowed(instr_allowed),
    .receipt_required(receipt_required),
    .current_mu_cost(mu_accumulator),
    .proposed_cost(proposed_cost),
    .partition_count(next_module_id),
    .memory_isolation(32'hCAFEBABE),  // Placeholder - would check actual memory isolation
    .receipt_value(receipt_value),
    .receipt_valid(receipt_valid),
    .receipt_accepted(receipt_accepted),
    .cost_gate_open(cost_gate_open),
    .partition_gate_open(partition_gate_open),
    .core_status(core_status),
    .enforcement_active(enforcement_active)
);

// Instantiate CLZ helper for 8-bit values (compute ceil(log2(x)) for x<=255)
wire [3:0] clz8_out;
reg [7:0] clz8_in;
clz8 clz8_inst (.x(clz8_in), .out(clz8_out));

// Deterministic helper for ceil(log2(x)) on small positive integers.
function automatic integer ceil_log2_8;
    input integer x;
    begin
        if (x <= 0) ceil_log2_8 = 1;
        else if (x <= 2) ceil_log2_8 = 1;
        else if (x <= 4) ceil_log2_8 = 2;
        else if (x <= 8) ceil_log2_8 = 3;
        else if (x <= 16) ceil_log2_8 = 4;
        else if (x <= 32) ceil_log2_8 = 5;
        else if (x <= 64) ceil_log2_8 = 6;
        else if (x <= 128) ceil_log2_8 = 7;
        else ceil_log2_8 = 8;
    end
endfunction

// Logic engine interface
assign logic_req = (state == STATE_LOGIC);
assign logic_addr = {24'h0, operand_a, operand_b};

// Python execution interface
assign py_req = (state == STATE_PYTHON);
assign py_code_addr = {24'h0, operand_a, operand_b};

// Memory interface (simplified)
assign mem_addr = pc_reg;
assign mem_wdata = 32'h0;
assign mem_we = 1'b0;
assign mem_en = 1'b1;

endmodule

// ---------------------------------------------------------------------------
// Local helper modules
// ---------------------------------------------------------------------------

// Simple combinational module returning ceiling(log2(x)) for up to 8-bit input
module clz8(
    input [7:0] x,
    output reg [3:0] out
);

always @(*) begin
    if (x == 0) out = 1;
    else if (x <= 1) out = 1;
    else if (x <= 2) out = 1;
    else if (x <= 4) out = 2;
    else if (x <= 8) out = 3;
    else if (x <= 16) out = 4;
    else if (x <= 32) out = 5;
    else if (x <= 64) out = 6;
    else if (x <= 128) out = 7;
    else out = 8;
end
endmodule