(* ================================================================= *)
(* Bridge module providing concrete implementations from archive    *)
(* This module extracts working definitions from the archive to     *)
(* avoid circular dependencies and compilation errors.              *)
(*                                                                   *)
(* STATUS: Partially complete                                        *)
(*   - Core definitions (run1, run_n, setup_state): CONCRETE ✓     *)
(*   - Basic lemmas (setup_state_regs_length, inv_min): PROVED ✓   *)
(*   - Helper lemmas (nth_add_skipn, nth_firstn_lt): PROVED ✓      *)
(*   - Transition lemmas: ADMITTED (require symbolic execution)     *)
(*                                                                   *)
(* NOTE: Relocated under thielemachine/verification to quarantine   *)
(* the instruction-level replay from the default `make core` flow.  *)
(* Use `make -C coq bridge` (or `verification`) to exercise this    *)
(* artifact without blocking the audited tier.                      *)
(*                                                                   *)
(* To complete: The transition lemmas require detailed symbolic     *)
(* execution proofs through the CPU interpreter. These are complex  *)
(* but mechanizable - they involve stepping through the instruction *)
(* sequence and maintaining invariants.                             *)
(* ================================================================= *)

From Coq Require Import List Arith Lia PeanoNat Bool ZArith String.
From ThieleUniversal Require Import TM UTM_Rules CPU UTM_Program UTM_Encode.
Import ListNotations.

Local Open Scope nat_scope.
Local Notation length := List.length.

(* Instrumentation helpers to locate long-running proofs during timed bridge
   builds.  The [Time] vernac modifier is applied to the key loop lemmas, and
   [bridge_checkpoint] marks entry into their proofs so a timed build can
   report the last completed milestone before hitting a timeout. *)
Ltac bridge_checkpoint msg :=
  let s := eval compute in msg in idtac "[bridge]" s.

(* ----------------------------------------------------------------- *)
(* Program encoding                                                  *)
(* ----------------------------------------------------------------- *)

(* The encoded universal program *)
Definition program : list nat :=
  flat_map UTM_Encode.encode_instr_words UTM_Program.program_instrs.

(* Compute the concrete program length once so decoding bounds can reuse it
   without re-running a large reduction. *)
Definition program_len : nat := Eval vm_compute in List.length program.

Lemma program_length_eq : List.length program = program_len.
Proof. reflexivity. Qed.

(* ----------------------------------------------------------------- *)
(* CPU Execution - from ThieleUniversal_Run1.v                      *)
(* ----------------------------------------------------------------- *)

(* Decode the instruction at the current program counter. *)
Definition decode_instr (st : CPU.State) : CPU.Instr :=
  UTM_Encode.decode_instr_from_mem st.(CPU.mem) (4 * CPU.read_reg CPU.REG_PC st).

(* Single step execution *)
Definition run1 (s : CPU.State) : CPU.State :=
  CPU.step (decode_instr s) s.

(* Multi-step execution *)
Fixpoint run_n (s : CPU.State) (n : nat) : CPU.State :=
  match n with
  | 0 => s
  | S n' => run_n (run1 s) n'
  end.

(* A reflection-friendly equality on states.  The CPU.State record contains
   only lists and naturals, so a structural Boolean equality lets us delegate
   large execution traces to [vm_compute]/[native_compute] without building a
   massive symbolic proof term. *)
Fixpoint list_eqb {A} (eqb : A -> A -> bool) (l1 l2 : list A) : bool :=
  match l1, l2 with
  | [], [] => true
  | x1 :: t1, x2 :: t2 => eqb x1 x2 && list_eqb eqb t1 t2
  | _, _ => false
  end.

Lemma list_eqb_spec {A} (eqb : A -> A -> bool) (eqb_spec : forall x y, eqb x y = true <-> x = y) :
  forall l1 l2, list_eqb eqb l1 l2 = true <-> l1 = l2.
Proof.
  induction l1 as [|x1 t1 IH]; destruct l2 as [|x2 t2]; simpl; try firstorder congruence.
  rewrite Bool.andb_true_iff, eqb_spec, IH. firstorder congruence.
Qed.

Lemma list_eqb_refl {A} (eqb : A -> A -> bool) (eqb_refl : forall x, eqb x x = true) :
  forall l, list_eqb eqb l l = true.
Proof.
  induction l as [|x t IH]; simpl; rewrite ?eqb_refl, ?IH; reflexivity.
Qed.

Definition state_eqb (s1 s2 : CPU.State) : bool :=
  Nat.eqb s1.(CPU.cost) s2.(CPU.cost)
    && list_eqb Nat.eqb s1.(CPU.regs) s2.(CPU.regs)
    && list_eqb Nat.eqb s1.(CPU.mem) s2.(CPU.mem).

Lemma state_eqb_refl : forall s, state_eqb s s = true.
Proof.
  intro s. destruct s as [r m c].
  simpl.
  apply Bool.andb_true_iff. split.
  - apply Bool.andb_true_iff. split.
    + apply Nat.eqb_refl.
    + apply list_eqb_refl. intros x. apply Nat.eqb_refl.
  - apply list_eqb_refl. intros x. apply Nat.eqb_refl.
Qed.

Lemma state_eqb_true_iff : forall s1 s2, state_eqb s1 s2 = true <-> s1 = s2.
Proof.
  intros s1 s2; split; intro H.
  - destruct s1 as [r1 m1 c1], s2 as [r2 m2 c2]; simpl in H.
    apply Bool.andb_true_iff in H as [Hcost_reg Hmem].
    apply Bool.andb_true_iff in Hcost_reg as [Hcost Hregs].
    apply Nat.eqb_eq in Hcost.
    apply (list_eqb_spec Nat.eqb Nat.eqb_eq) in Hregs.
    apply (list_eqb_spec Nat.eqb Nat.eqb_eq) in Hmem.
    simpl in Hcost, Hregs, Hmem.
    subst c2 r2 m2. reflexivity.
  - rewrite H. destruct s2 as [r m c].
    apply state_eqb_refl.
  Qed.

Definition check_transition (start_state end_state : CPU.State) (steps : nat) : bool :=
  state_eqb (run_n start_state steps) end_state.

Lemma check_transition_sound : forall s1 s2 n,
  check_transition s1 s2 n = true -> run_n s1 n = s2.
Proof.
  unfold check_transition.
  intros s1 s2 n H.
  apply state_eqb_true_iff in H; assumption.
Qed.

Ltac vm_run_n :=
  match goal with
  | |- run_n ?s ?n = ?t =>
      apply (check_transition_sound s t n);
      vm_compute; reflexivity
  end.

(* Symbolic steppers for small, concrete prefixes.  These avoid the
   `vm_compute`/`native_compute` path when the starting state is still
   symbolic, but the program being fetched is concrete. *)
Ltac step_symbolic :=
  cbv [run1 CPU.step UTM_Encode.decode_instr_from_mem] in *;
  simpl.

(* ----------------------------------------------------------------- *)
(* State Setup - extracted from ThieleUniversal.v                   *)
(* ----------------------------------------------------------------- *)

(* Helper: set nth element of a list *)
Definition set_nth {A : Type} (l : list A) (n : nat) (v : A) : list A :=
  firstn n l ++ [v] ++ skipn (S n) l.

(* Helper: pad list to length n with zeros *)
Definition pad_to (n : nat) (l : list nat) : list nat :=
  l ++ repeat 0 (n - length l).

Lemma pad_to_expand : forall n l,
  pad_to n l = l ++ repeat 0 (n - length l).
Proof. reflexivity. Qed.

Lemma length_pad_to_ge : forall l n,
  length l <= n -> length (pad_to n l) = n.
Proof.
  intros l n Hle.
  unfold pad_to.
  rewrite app_length, repeat_length.
  lia.
Qed.

Lemma length_pad_to_ge_base : forall l n,
  length (pad_to n l) >= length l.
Proof.
  intros l n.
  unfold pad_to.
  rewrite app_length, repeat_length.
  lia.
Qed.

Lemma nth_app_lt : forall {A} (l1 l2 : list A) n d,
  n < length l1 -> nth n (l1 ++ l2) d = nth n l1 d.
Proof.
  intros A l1 l2 n d Hlt.
  revert n Hlt.
  induction l1 as [|x l1 IH]; intros [|n] Hlt; simpl in *; try lia; auto.
  apply IH. lia.
Qed.

Lemma firstn_pad_to : forall l n,
  length l <= n -> firstn (length l) (pad_to n l) = l.
Proof.
  intros l n Hle.
  unfold pad_to.
  rewrite firstn_app.
  rewrite Nat.sub_diag.
  simpl.
  rewrite firstn_all.
  rewrite app_nil_r.
  reflexivity.
Qed.

Lemma firstn_app_le' : forall {A} n (l1 l2 : list A),
  n <= length l1 -> firstn n (l1 ++ l2) = firstn n l1.
Proof.
  intros A n l1 l2 Hn.
  rewrite firstn_app.
  replace (n - length l1) with 0 by lia.
  simpl.
  rewrite app_nil_r.
  reflexivity.
Qed.

Lemma skipn_app_le' : forall {A} n (l1 l2 : list A),
  n <= length l1 -> skipn n (l1 ++ l2) = skipn n l1 ++ l2.
Proof.
  intros A n l1 l2 Hn.
  rewrite skipn_app.
  replace (n - length l1) with 0 by lia.
  simpl.
  reflexivity.
Qed.

Lemma firstn_pad_to_le : forall l n k,
  k <= length l -> firstn k (pad_to n l) = firstn k l.
Proof.
  intros l n k Hk.
  unfold pad_to.
  rewrite firstn_app_le' by lia.
  reflexivity.
Qed.

Lemma firstn_pad_to_app_le : forall l n rest k,
  k <= length l -> firstn k (pad_to n l ++ rest) = firstn k l.
Proof.
  intros l n rest k Hk.
  unfold pad_to.
  rewrite firstn_app_le' by (rewrite app_length, repeat_length; lia).
  rewrite firstn_app_le' by lia.
  reflexivity.
Qed.

Lemma skipn_pad_to_app : forall l n rest,
  length l <= n -> skipn n (pad_to n l ++ rest) = rest.
Proof.
  intros l n rest Hle.
  unfold pad_to.
  rewrite skipn_app.
  assert (Hlen : length (l ++ repeat 0 (n - length l)) = n).
  { rewrite app_length, repeat_length. lia. }
  rewrite Hlen.
  rewrite Nat.sub_diag.
  rewrite skipn_all2 by lia.
  reflexivity.
Qed.

Lemma firstn_program_prefix :
  length program <= UTM_Program.RULES_START_ADDR ->
  forall rules,
    firstn (length program)
      (pad_to UTM_Program.TAPE_START_ADDR
         (pad_to UTM_Program.RULES_START_ADDR program ++ rules)) = program.
Proof.
  intros Hprog rules.
  remember (length program) as len_prog eqn:Hlen_prog.
  assert (Hprog_len : length program <= UTM_Program.RULES_START_ADDR)
    by (rewrite <- Hlen_prog; exact Hprog).
  assert (Hpad_window : firstn len_prog
           (pad_to UTM_Program.TAPE_START_ADDR
              (pad_to UTM_Program.RULES_START_ADDR program ++ rules)) =
          firstn len_prog (pad_to UTM_Program.RULES_START_ADDR program ++ rules)).
  { apply firstn_pad_to_le.
    rewrite app_length, length_pad_to_ge with (l := program)
        (n := UTM_Program.RULES_START_ADDR) by exact Hprog_len.
    rewrite Hlen_prog. lia. }
  assert (Hmem_prog : firstn len_prog
            (pad_to UTM_Program.RULES_START_ADDR program ++ rules) =
          firstn len_prog program).
  { rewrite firstn_pad_to_app_le with (l := program)
        (n := UTM_Program.RULES_START_ADDR) (rest := rules) (k := len_prog)
      by (rewrite Hlen_prog; lia).
    reflexivity. }
  assert (Hfirstn_prog : firstn len_prog program = program).
  { rewrite Hlen_prog. apply firstn_all. }
  eapply eq_trans. exact Hpad_window.
  eapply eq_trans. exact Hmem_prog.
  exact Hfirstn_prog.
Qed.

Lemma firstn_skipn_pad_to_app : forall l n rest,
  length l <= n -> firstn (length rest) (skipn n (pad_to n l ++ rest)) = rest.
Proof.
  intros l n rest Hle.
  rewrite skipn_pad_to_app by assumption.
  apply firstn_all.
Qed.

Lemma skipn_pad_to_split : forall l n k,
  k <= length l ->
  skipn k (pad_to n l) = skipn k l ++ repeat 0 (n - length l).
Proof.
  intros l n k Hk.
  unfold pad_to.
  rewrite skipn_app_le' by lia.
  reflexivity.
Qed.

Lemma firstn_rules_window :
  length program <= UTM_Program.RULES_START_ADDR ->
  forall rules,
    length rules <= UTM_Program.TAPE_START_ADDR - UTM_Program.RULES_START_ADDR ->
    firstn (length rules)
      (skipn UTM_Program.RULES_START_ADDR
         (pad_to UTM_Program.TAPE_START_ADDR
            (pad_to UTM_Program.RULES_START_ADDR program ++ rules))) = rules.
Proof.
  intros Hprog rules Hfit.
  set (memprog := pad_to UTM_Program.RULES_START_ADDR program).
  set (memrules := memprog ++ rules).
  assert (Hmemprog_len : length memprog = UTM_Program.RULES_START_ADDR).
  { subst memprog. apply length_pad_to_ge. exact Hprog. }
  assert (Hskip_memrules : skipn UTM_Program.RULES_START_ADDR memrules = rules).
  { unfold memrules.
    rewrite skipn_app_le' by (rewrite Hmemprog_len; lia).
    rewrite <- Hmemprog_len.
    rewrite skipn_all.
    simpl. reflexivity. }
  assert (Hskip_pad :
    skipn UTM_Program.RULES_START_ADDR
      (pad_to UTM_Program.TAPE_START_ADDR memrules) =
    skipn UTM_Program.RULES_START_ADDR memrules ++
      repeat 0 (UTM_Program.TAPE_START_ADDR - length memrules)).
  { apply skipn_pad_to_split.
    unfold memrules.
    rewrite app_length, Hmemprog_len.
    lia. }
  rewrite Hskip_pad.
  rewrite Hskip_memrules.
  rewrite firstn_app_le' by lia.
  apply firstn_all.
Qed.

Lemma firstn_skipn_app_exact : forall {A} (pref rest : list A) n,
  length pref = n ->
  firstn (length rest) (skipn n (pref ++ rest)) = rest.
Proof.
  intros A pref rest n Hlen.
  rewrite skipn_app.
  rewrite Hlen.
  rewrite Nat.sub_diag.
  rewrite <- Hlen.
  rewrite skipn_all.
  simpl.
  apply firstn_all.
Qed.

(* Padding preserves existing elements below the original length. *)
Lemma nth_pad_to_lt : forall (l : list nat) n d k,
  n < length l ->
  nth n (pad_to k l) d = nth n l d.
Proof.
  intros l n d k Hlt.
  unfold pad_to.
  apply nth_app_lt; lia.
Qed.

(* Avoid expanding large padded memories during later proofs. *)
#[local] Opaque pad_to repeat.

(* Setup initial CPU state from TM configuration *)
Definition setup_state (tm : TM) (conf : TMConfig) : CPU.State :=
  let '((q, tape), head) := conf in
  let regs0 := repeat 0 10 in
  let regs1 := set_nth regs0 CPU.REG_Q q in
  let regs2 := set_nth regs1 CPU.REG_HEAD head in
  let regs3 := set_nth regs2 CPU.REG_PC 0 in
  let rules := UTM_Encode.encode_rules tm.(tm_rules) in
  let mem0 := pad_to UTM_Program.RULES_START_ADDR program in
  let mem1 := pad_to UTM_Program.TAPE_START_ADDR (mem0 ++ rules) in
  {| CPU.regs := regs3; CPU.mem := mem1 ++ tape; CPU.cost := 0 |}.

(* Don't make these opaque yet - we need them for foundational lemmas *)

(* ----------------------------------------------------------------- *)
(* Program layout shortcuts                                          *)
(* ----------------------------------------------------------------- *)

(* Tactic to discharge fixed program-length bounds when decoding. *)
Ltac calc_bounds :=
  rewrite program_length_eq;
  unfold program_len;
  simpl;
  lia.

(* The concrete program lives at the front of memory; when the PC stays within
   the program bounds we can read directly from the static [program] list and
   ignore the symbolic rules/tape suffix. *)
Lemma program_memory_lookup : forall tm conf n,
  n < length program ->
  nth n (CPU.mem (setup_state tm conf)) 0 = nth n program 0.
Proof.
  intros tm conf n Hn.
  destruct conf as ((q, tape), head).
  unfold setup_state; simpl.
  set (rules := UTM_Encode.encode_rules tm.(tm_rules)).
  set (mem0 := pad_to UTM_Program.RULES_START_ADDR program).
  set (mem1 := pad_to UTM_Program.TAPE_START_ADDR (mem0 ++ rules)).
  assert (Hmem0_len : n < length mem0).
  { subst mem0. eapply Nat.lt_le_trans; [exact Hn|]. apply length_pad_to_ge_base. }
  assert (Hmem1_len : n < length mem1).
  { subst mem1.
    eapply Nat.lt_le_trans; [| apply length_pad_to_ge_base ].
    eapply Nat.lt_le_trans; [exact Hmem0_len|].
    rewrite app_length; lia.
  }
  subst mem1.
  eapply eq_trans.
  { apply (@nth_app_lt nat (pad_to UTM_Program.TAPE_START_ADDR (mem0 ++ rules)) tape n 0).
    exact Hmem1_len. }
  eapply eq_trans.
  { apply (nth_pad_to_lt (mem0 ++ rules) n 0 UTM_Program.TAPE_START_ADDR).
    rewrite app_length. lia. }
  rewrite nth_app_lt by lia.
  subst mem0.
  rewrite (nth_pad_to_lt program n 0 UTM_Program.RULES_START_ADDR) by exact Hn.
  reflexivity.
Qed.

(* If a state already exposes the concrete program prefix, we can reuse that
   fact to read directly from [program] without re-running the padding
   expansions.  This lets later steps avoid reopening [setup_state]. *)

Lemma decode_program_at_pc : forall tm conf pc,
  4 * pc + 3 < length program ->
  UTM_Encode.decode_instr_from_mem (CPU.mem (setup_state tm conf)) (4 * pc) =
  UTM_Encode.decode_instr_from_mem program (4 * pc).
Proof.
  intros tm conf pc Hbound.
  unfold UTM_Encode.decode_instr_from_mem.
  repeat rewrite program_memory_lookup; try lia.
  reflexivity.
Qed.

(* ----------------------------------------------------------------- *)
(* Basic lemmas about setup_state                                    *)
(* ----------------------------------------------------------------- *)

Lemma length_set_nth : forall {A : Type} (l : list A) n v,
  n < length l ->
  length (set_nth l n v) = length l.
Proof.
  intros A l n v Hn.
  unfold set_nth.
  rewrite app_length, app_length.
  rewrite firstn_length, skipn_length.
  simpl.
  rewrite Nat.min_l by lia.
  lia.
Qed.

Lemma setup_state_regs_length :
  forall tm conf, length (CPU.regs (setup_state tm conf)) = 10.
Proof.
  intros tm conf.
  destruct conf as ((q, tape), head).
  unfold setup_state. simpl CPU.regs.
  repeat (rewrite length_set_nth; [|repeat rewrite length_set_nth; simpl; lia]).
  simpl. reflexivity.
Qed.

(* ----------------------------------------------------------------- *)
(* State predicates and invariants                                   *)
(* ----------------------------------------------------------------- *)

Definition inv_min (st : CPU.State) (tm : TM) (conf : TMConfig) : Prop :=
  let '(q, tape, head) := conf in
  CPU.read_reg CPU.REG_Q st = q /\
  CPU.read_reg CPU.REG_HEAD st = head.

Lemma inv_min_setup_state : forall tm conf,
  inv_min (setup_state tm conf) tm conf.
Proof.
  intros tm ((q, tape), head).
  unfold inv_min, setup_state; simpl.
  split; unfold CPU.read_reg; repeat (rewrite nth_skipn || simpl); try lia; reflexivity.
Qed.

Definition IS_FetchSymbol (pc : nat) : Prop := pc = 0.
Definition IS_FindRule_Start (pc : nat) : Prop := pc = 3.

(* Tape window predicate: memory correctly encodes the tape *)
Definition tape_window_ok (st : CPU.State) (tape : list nat) : Prop :=
  firstn (length tape) (skipn UTM_Program.TAPE_START_ADDR st.(CPU.mem)) = tape.

Lemma tape_window_ok_setup_state : forall tm q tape head,
  length program <= UTM_Program.RULES_START_ADDR ->
  length (UTM_Encode.encode_rules tm.(tm_rules))
    <= UTM_Program.TAPE_START_ADDR - UTM_Program.RULES_START_ADDR ->
  tape_window_ok (setup_state tm ((q, tape), head)) tape.
Proof.
  intros tm q tape head Hprog Hrules.
  unfold tape_window_ok, setup_state.
  set (rrules := UTM_Encode.encode_rules tm.(tm_rules)).
  set (mem0 := pad_to UTM_Program.RULES_START_ADDR program).
  set (mem1 := pad_to UTM_Program.TAPE_START_ADDR (mem0 ++ rrules)).
  simpl.
  assert (Hmem0_len : length mem0 = UTM_Program.RULES_START_ADDR).
  { subst mem0. apply length_pad_to_ge. exact Hprog. }
  assert (Hfit : length (mem0 ++ rrules) <= UTM_Program.TAPE_START_ADDR).
  { rewrite app_length, Hmem0_len.
    pose proof UTM_Program.RULES_START_ADDR_le_TAPE_START_ADDR as Hle.
    rewrite <- (Arith_prebase.le_plus_minus_r_stt _ _ Hle).
    apply Nat.add_le_mono_l. exact Hrules. }
  subst mem1.
  assert (Hmem1_len : length (pad_to UTM_Program.TAPE_START_ADDR (mem0 ++ rrules))
                        = UTM_Program.TAPE_START_ADDR).
  { apply length_pad_to_ge. exact Hfit. }
  apply (@firstn_skipn_app_exact
           nat
           (pad_to UTM_Program.TAPE_START_ADDR (mem0 ++ rrules))
           tape
           UTM_Program.TAPE_START_ADDR).
  exact Hmem1_len.
Qed.

(* Full invariant relating CPU state to TM configuration *)
Definition inv (st : CPU.State) (tm : TM) (conf : TMConfig) : Prop :=
  let '((q, tape), head) := conf in
  CPU.read_reg CPU.REG_Q st = q /\
  CPU.read_reg CPU.REG_HEAD st = head /\
  CPU.read_reg CPU.REG_PC st = 0 /\
  tape_window_ok st tape /\
  firstn (length program) st.(CPU.mem) = program /\
  firstn (length (UTM_Encode.encode_rules tm.(tm_rules)))
         (skipn UTM_Program.RULES_START_ADDR st.(CPU.mem)) = 
    UTM_Encode.encode_rules tm.(tm_rules).

Lemma inv_setup_state : forall tm conf,
  length program <= UTM_Program.RULES_START_ADDR ->
  length (UTM_Encode.encode_rules tm.(tm_rules))
    <= UTM_Program.TAPE_START_ADDR - UTM_Program.RULES_START_ADDR ->
  inv (setup_state tm conf) tm conf.
Proof.
  intros tm ((q, tape), head) Hprog Hrules.
  pose proof (inv_min_setup_state tm ((q, tape), head)) as Hmin.
  destruct Hmin as [Hq Hhead].
  unfold inv.
  simpl.
  split. exact Hq.
  split. exact Hhead.
  split.
  { unfold setup_state.
    simpl.
    unfold CPU.read_reg.
    repeat (rewrite nth_skipn || simpl); try lia; reflexivity. }
  split. apply tape_window_ok_setup_state; assumption.
  split.
  - unfold setup_state; simpl.
    set (rules := UTM_Encode.encode_rules tm.(tm_rules)).
    set (mem0 := pad_to UTM_Program.RULES_START_ADDR program).
    assert (Hmem0_len : length mem0 = UTM_Program.RULES_START_ADDR)
      by (subst mem0; apply length_pad_to_ge; exact Hprog).
    assert (Hfit : length (mem0 ++ rules) <= UTM_Program.TAPE_START_ADDR).
    { rewrite app_length, Hmem0_len.
      assert (Heq : UTM_Program.TAPE_START_ADDR =
        UTM_Program.RULES_START_ADDR + (UTM_Program.TAPE_START_ADDR - UTM_Program.RULES_START_ADDR))
        by (unfold UTM_Program.TAPE_START_ADDR, UTM_Program.RULES_START_ADDR; lia).
      rewrite Heq. apply Nat.add_le_mono_l. exact Hrules. }
    assert (Hmem1_len : length (pad_to UTM_Program.TAPE_START_ADDR (mem0 ++ rules))
                        = UTM_Program.TAPE_START_ADDR)
      by (apply length_pad_to_ge; exact Hfit).
    assert (Hprefix :
      firstn (length program)
        ((pad_to UTM_Program.TAPE_START_ADDR (mem0 ++ rules)) ++ tape)
      = firstn (length program)
          (pad_to UTM_Program.TAPE_START_ADDR (mem0 ++ rules)))
      by (apply firstn_app_le'; rewrite Hmem1_len;
          apply (Nat.le_trans _ _ _ Hprog); exact UTM_Program.RULES_START_ADDR_le_TAPE_START_ADDR).
    eapply eq_trans; [exact Hprefix|].
    subst mem0. apply (firstn_program_prefix Hprog rules).
  - unfold setup_state; simpl.
    set (rules := UTM_Encode.encode_rules tm.(tm_rules)).
    set (mem0 := pad_to UTM_Program.RULES_START_ADDR program).
    assert (Hmem0_len : length mem0 = UTM_Program.RULES_START_ADDR)
      by (subst mem0; apply length_pad_to_ge; exact Hprog).
    assert (Hfit : length (mem0 ++ rules) <= UTM_Program.TAPE_START_ADDR).
    { rewrite app_length, Hmem0_len.
      assert (Heq : UTM_Program.TAPE_START_ADDR =
        UTM_Program.RULES_START_ADDR + (UTM_Program.TAPE_START_ADDR - UTM_Program.RULES_START_ADDR))
        by (unfold UTM_Program.TAPE_START_ADDR, UTM_Program.RULES_START_ADDR; lia).
      rewrite Heq. apply Nat.add_le_mono_l. exact Hrules. }
    assert (Hmem1_len : length (pad_to UTM_Program.TAPE_START_ADDR (mem0 ++ rules))
                        = UTM_Program.TAPE_START_ADDR)
      by (apply length_pad_to_ge; exact Hfit).
    assert (Hskip :
      skipn UTM_Program.RULES_START_ADDR
        ((pad_to UTM_Program.TAPE_START_ADDR (mem0 ++ rules)) ++ tape)
      = skipn UTM_Program.RULES_START_ADDR
          (pad_to UTM_Program.TAPE_START_ADDR (mem0 ++ rules)) ++ tape)
      by (apply skipn_app_le'; rewrite Hmem1_len; exact UTM_Program.RULES_START_ADDR_le_TAPE_START_ADDR).
    assert (Hskip_first :
      firstn (length rules)
        (skipn UTM_Program.RULES_START_ADDR
                 ((pad_to UTM_Program.TAPE_START_ADDR (mem0 ++ rules)) ++ tape))
      = firstn (length rules)
          (skipn UTM_Program.RULES_START_ADDR
                   (pad_to UTM_Program.TAPE_START_ADDR (mem0 ++ rules)) ++ tape))
      by (rewrite Hskip; reflexivity).
    assert (Hdrop :
      firstn (length rules)
        (skipn UTM_Program.RULES_START_ADDR
                 (pad_to UTM_Program.TAPE_START_ADDR (mem0 ++ rules)) ++ tape)
      = firstn (length rules)
          (skipn UTM_Program.RULES_START_ADDR
                 (pad_to UTM_Program.TAPE_START_ADDR (mem0 ++ rules))))
      by (apply firstn_app_le'; rewrite skipn_length, Hmem1_len;
          apply (Nat.le_trans _ _ _ Hrules); lia).
    eapply eq_trans; [exact Hskip_first|].
    eapply eq_trans; [exact Hdrop|].
    subst mem0. apply (firstn_rules_window Hprog rules). exact Hrules.
Qed.

Definition inv_core (st : CPU.State) (tm : TM) (conf : TMConfig) : Prop :=
  let '((q, tape), head) := conf in
  CPU.read_reg CPU.REG_Q st = q /\
  CPU.read_reg CPU.REG_HEAD st = head /\
  tape_window_ok st tape /\
  firstn (length program) st.(CPU.mem) = program /\
  firstn (length (UTM_Encode.encode_rules tm.(tm_rules)))
        (skipn UTM_Program.RULES_START_ADDR st.(CPU.mem)) =
    UTM_Encode.encode_rules tm.(tm_rules) /\
  length (skipn UTM_Program.TAPE_START_ADDR st.(CPU.mem)) = length tape.

Definition find_rule_start_inv (tm : TM) (conf : TMConfig) (cpu : CPU.State) : Prop :=
  IS_FindRule_Start (CPU.read_reg CPU.REG_PC cpu) /\
  inv_min cpu tm conf.

(* Specialised small-stepper for states whose memory prefix is the encoded
   program.  When explicit decoder hypotheses are available, rewrite with them
   instead of unfolding the program prefix; this keeps small goal states during
   timed builds. *)
Ltac step_fast :=
  unfold run1, CPU.step;
  (* Prefer explicit decoder hypotheses over unfolding the concrete program, so
     small symbolic goals avoid expensive [calc_bounds] calls. *)
  first
    [ match goal with
      | H : decode_instr ?s = _ |- context [decode_instr ?s] => rewrite H
      end
    (* If no hypothesis is available, compute the decoder result directly
       instead of triggering [calc_bounds] on the program prefix.  This keeps
       timed bridge builds from spending most of their budget in the fallback
       bound solver when stepping through short concrete traces. *)
    | lazymatch goal with
      | |- context [decode_instr ?s] =>
          let inst := eval vm_compute in (decode_instr s) in
          change (decode_instr s) with inst
      end
    | try rewrite decode_program_at_pc by calc_bounds ];
  cbn [CPU.read_reg CPU.mem CPU.regs CPU.cost];
  simpl.

Ltac step_n n :=
  lazymatch n with
  | 0 => cbn [run_n] in *
  | S ?n' =>
      cbn [run_n] in *;
      step_fast;
      step_n n'
  end.

Lemma run1_decode : forall st,
  run1 st = CPU.step (decode_instr st) st.
Proof.
  intro st.
  unfold run1, decode_instr.
  reflexivity.
Qed.

(* ----------------------------------------------------------------- *)
(* Helper lemmas                                                      *)
(* ----------------------------------------------------------------- *)

Lemma nth_add_skipn : forall {A} n m (l : list A) d,
  nth n (skipn m l) d = nth (m + n) l d.
Proof.
  intros A n m l d.
  revert n m.
  induction l as [|x l IH]; intros n m.
  - destruct m; destruct n; simpl; reflexivity.
  - destruct m.
    + simpl. reflexivity.
    + simpl. apply IH.
Qed.

Lemma nth_firstn_lt : forall {A} n m (l : list A) d,
  n < m -> nth n (firstn m l) d = nth n l d.
Proof.
  intros A n m l d Hn.
  revert n m Hn.
  induction l as [|x l IH]; intros n m Hn.
  - destruct n; destruct m; simpl; try reflexivity; try lia.
  - destruct n; destruct m; simpl; try reflexivity; try lia.
    apply IH. lia.
Qed.

(* Placeholder transition lemmas - these would need full proofs *)
(* For now we provide stubs that can be filled in *)

(* ----------------------------------------------------------------- *)
(* Common Infrastructure Lemmas                                      *)
(* ----------------------------------------------------------------- *)

(* Step composition lemmas *)
Lemma run_n_add : forall cpu m n,
  run_n cpu (m + n) = run_n (run_n cpu m) n.
Proof.
  intros cpu m n.
  revert cpu.
  induction m as [|m' IH]; intros cpu.
  - simpl. reflexivity.
  - simpl. rewrite IH. reflexivity.
Qed.

Lemma run_n_S : forall cpu n,
  run_n cpu (S n) = run_n (run1 cpu) n.
Proof.
  intros cpu n.
  simpl. reflexivity.
Qed.

Lemma run_n_0 : forall cpu,
  run_n cpu 0 = cpu.
Proof.
  intros cpu. reflexivity.
Qed.

Lemma run_n_1 : forall cpu,
  run_n cpu 1 = run1 cpu.
Proof.
  intros cpu. reflexivity.
Qed.

(* Prevent large proof terms from repeatedly unfolding the small-step
   interpreter.  The structural lemmas above expose the only rewrites we
   rely on, so the operational definitions can remain opaque during the
   heavy FindRule proofs. *)
#[local] Opaque run_n decode_instr.

(* Make key definitions opaque to prevent expensive unfolding during proofs.
   This stops the unifier from expanding massive symbolic lists. *)
#[global] Opaque program.
#[global] Opaque pad_to.
#[global] Opaque setup_state.

(* Rewrite run_n in terms of iterations *)
Lemma run_n_unfold_3 : forall cpu,
  run_n cpu 3 = run1 (run1 (run1 cpu)).
Proof.
  intros cpu.
  simpl. reflexivity.
Qed.

(* Memory and register helpers *)
Lemma read_reg_bounds : forall cpu r,
  r < 10 ->
  exists v, CPU.read_reg r cpu = v.
Proof.
  intros cpu r Hr.
  exists (CPU.read_reg r cpu).
  reflexivity.
Qed.

(* Key lemma: reading from the register you just wrote gives the value *)
Lemma read_reg_write_reg_same : forall r v st,
  r < length st.(CPU.regs) ->
  CPU.read_reg r (CPU.write_reg r v st) = v.
Proof.
  intros r v st Hr.
  unfold CPU.read_reg, CPU.write_reg. simpl.
  (* After write_reg r v, the register file is: firstn r regs ++ [v] ++ skipn (S r) regs *)
  (* Reading at position r gives v *)
  rewrite app_nth2.
  - rewrite firstn_length.
    rewrite Nat.min_l by lia.
    replace (r - r) with 0 by lia.
    simpl. reflexivity.
  - rewrite firstn_length.
    rewrite Nat.min_l by lia.
    lia.
Qed.

(* Reading a different register after write *)
Lemma read_reg_write_reg_diff : forall r1 r2 v st,
  r1 <> r2 ->
  r1 < length st.(CPU.regs) ->
  r2 < length st.(CPU.regs) ->
  CPU.read_reg r1 (CPU.write_reg r2 v st) = CPU.read_reg r1 st.
Proof.
  intros r1 r2 v st Hneq Hr1 Hr2.
  unfold CPU.read_reg, CPU.write_reg. simpl.
  (* Need to show: nth r1 (firstn r2 regs ++ [v] ++ skipn (S r2) regs) 0 = nth r1 regs 0 *)
  destruct (Nat.ltb r1 r2) eqn:Hlt.
  - (* Case r1 < r2: r1 is in the firstn part *)
    apply Nat.ltb_lt in Hlt.
    rewrite app_nth1.
    + apply nth_firstn_lt. exact Hlt.
    + rewrite firstn_length. rewrite Nat.min_l; [lia|lia].
  - (* Case r1 >= r2, but r1 <> r2, so r1 > r2 *)
    apply Nat.ltb_nlt in Hlt.
    assert (r1 > r2) by lia.
    (* r1 is beyond the firstn r2 part *)
    rewrite app_nth2.
    + rewrite firstn_length. rewrite Nat.min_l; [|lia].
      (* nth (r1 - r2) ([v] ++ skipn (S r2) regs) 0 = nth r1 regs 0 *)
      destruct (r1 - r2) as [|n] eqn:Hdiff; [lia|].
      simpl.
      (* nth n (skipn (S r2) regs) 0 = nth r1 regs 0 *)
      assert (Heqr1: r1 = S r2 + n) by lia.
      rewrite Heqr1.
      (* Now prove: nth n (skipn (S r2) regs) 0 = nth (S r2 + n) regs 0 *)
      clear Heqr1 Hdiff Hneq Hr1 Hr2 H Hlt v r1.
      generalize dependent n. generalize dependent r2.
      induction (CPU.regs st) as [|x xs IH]; intros.
      { destruct n, r2; reflexivity. }
      destruct r2; simpl.
      { destruct n; reflexivity. }
      { apply IH. }
    + rewrite firstn_length. rewrite Nat.min_l; [lia|lia].
Qed.

(*Writing to a register never shrinks the register file. *)
Lemma length_write_reg_ge : forall r v st,
  length (CPU.write_reg r v st).(CPU.regs) >= length st.(CPU.regs).
Proof.
  intros r v st.
  unfold CPU.write_reg. simpl.
  (* After unfolding: firstn r (CPU.regs st) ++ [v] ++ skipn (S r) (CPU.regs st) *)
  set (regs := CPU.regs st).
  assert (Hlen: forall (l : list nat) n m,
    length (firstn n l ++ m :: skipn (S n) l) >= length l).
  { intros l. induction l as [|x xs IHxs]; intros n m.
    - destruct n; simpl; lia.
    - destruct n; simpl.
      + lia.
      + simpl in IHxs. specialize (IHxs n m). simpl. lia. }
  apply (Hlen regs r v).
Qed.

(* Stepping cannot shorten the register file. *)
Lemma length_step_ge : forall instr st,
  length (CPU.regs (CPU.step instr st)) >= length st.(CPU.regs).
Proof.
  intros instr st.
  unfold CPU.step.
  remember (CPU.write_reg CPU.REG_PC (S (CPU.read_reg CPU.REG_PC st)) st) as st_pc eqn:Heq_st_pc.
  assert (Hlen_pc : length (CPU.regs st_pc) >= length st.(CPU.regs)).
  { subst st_pc. apply length_write_reg_ge. }
  clear Heq_st_pc.
  destruct instr; simpl.
  - (* LoadConst *) eapply Nat.le_trans; [apply Hlen_pc|apply length_write_reg_ge].
  - (* LoadIndirect *) eapply Nat.le_trans; [apply Hlen_pc|apply length_write_reg_ge].
  - (* StoreIndirect *) unfold CPU.write_mem; simpl; assumption.
  - (* CopyReg *) eapply Nat.le_trans; [apply Hlen_pc|apply length_write_reg_ge].
  - (* AddConst *) eapply Nat.le_trans; [apply Hlen_pc|apply length_write_reg_ge].
  - (* AddReg *) eapply Nat.le_trans; [apply Hlen_pc|apply length_write_reg_ge].
  - (* SubReg *) eapply Nat.le_trans; [apply Hlen_pc|apply length_write_reg_ge].
  - (* Jz: if zero, write_reg to st; otherwise st_pc *)
    destruct (Nat.eqb (CPU.read_reg rc st) 0).
    + apply length_write_reg_ge.
    + assumption.
  - (* Jnz: if zero, st_pc; otherwise write_reg to st *)
    destruct (Nat.eqb (CPU.read_reg rc st) 0).
    + assumption.
    + apply length_write_reg_ge.
  - (* Halt: returns st unchanged *)
    apply Nat.le_refl.
Qed.

(* Multi-step execution preserves or grows the register file length. *)
Lemma length_run_n_ge : forall st n,
  length (CPU.regs (run_n st n)) >= length st.(CPU.regs).
Proof.
  intros st n.
  revert st. (* Generalize st before induction so IH is universal *)
  induction n as [|n' IHn]; intros st.
  - (* Base case: n = 0 *)
    simpl. apply Nat.le_refl.
  - (* Inductive case: n = S n' *)
    simpl. (* run_n st (S n') = run_n (run1 st) n' *)
    (* IHn : forall st', length (run_n st' n') >= length st' *)
    (* Need: length (run_n (run1 st) n') >= length st *)
    assert (H1: length (CPU.regs (run1 st)) >= length (CPU.regs st)).
    { unfold run1. apply length_step_ge. }
    assert (H2: length (CPU.regs (run_n (run1 st) n')) >= length (CPU.regs (run1 st))).
    { apply IHn. }
    eapply Nat.le_trans; [exact H1 | exact H2].
Qed.

(* Helper: length is preserved by write_reg *)
Lemma length_write_reg : forall r v st,
  r < length st.(CPU.regs) ->
  length (CPU.write_reg r v st).(CPU.regs) = length st.(CPU.regs).
Proof.
  intros r v st Hr.
  unfold CPU.write_reg. simpl.
  (* Directly compute the length *)
  generalize dependent r. generalize dependent v.
  induction (CPU.regs st) as [|x xs IH]; intros.
  - simpl in Hr. lia.
  - destruct r; simpl.
    + simpl. reflexivity.
    + simpl. rewrite IH by (simpl in Hr; lia). reflexivity.
Qed.

(* CPU.step PC progression for non-branching instructions *)
(* Note: This lemma requires that rd <> REG_PC for all register-writing instructions.
   This is a constraint on the instruction encoding that should be enforced by the
   instruction decoder or compiler. The UTM program in UTM_Program.v satisfies this. *)
Lemma step_pc_increment : forall cpu instr,
  CPU.pc_unchanged instr ->
  CPU.read_reg CPU.REG_PC (CPU.step instr cpu) = S (CPU.read_reg CPU.REG_PC cpu).
Proof.
  intros cpu instr Hpc_unch.
  apply CPU.step_pc_succ.
  exact Hpc_unch.
Qed.

(* ----------------------------------------------------------------- *)
(* Instruction Decoding Lemmas                                       *)
(* ----------------------------------------------------------------- *)

(* Import the actual UTM program from archive *)
(* The program starts at PC=0 with these instructions:
   PC=0: LoadConst REG_TEMP1 TAPE_START_ADDR  (Fetch phase)
   PC=1: AddReg REG_ADDR REG_TEMP1 REG_HEAD
   PC=2: LoadIndirect REG_SYM REG_ADDR
   PC=3: LoadConst REG_ADDR RULES_START_ADDR  (FindRule phase starts)
   ...
*)

(* Lemmas about what instructions are at specific PCs *)
Lemma instr_at_pc_0 : 
  nth 0 UTM_Program.program_instrs CPU.Halt = 
  CPU.LoadConst CPU.REG_TEMP1 UTM_Program.TAPE_START_ADDR.
Proof.
  unfold UTM_Program.program_instrs. simpl. reflexivity.
Qed.

Lemma instr_at_pc_1 :
  nth 1 UTM_Program.program_instrs CPU.Halt =
  CPU.AddReg CPU.REG_ADDR CPU.REG_TEMP1 CPU.REG_HEAD.
Proof.
  unfold UTM_Program.program_instrs. simpl. reflexivity.
Qed.

Lemma instr_at_pc_2 :
  nth 2 UTM_Program.program_instrs CPU.Halt =
  CPU.LoadIndirect CPU.REG_SYM CPU.REG_ADDR.
Proof.
  unfold UTM_Program.program_instrs. simpl. reflexivity.
Qed.

Lemma instr_at_pc_3 :
  nth 3 UTM_Program.program_instrs CPU.Halt =
  CPU.LoadConst CPU.REG_ADDR UTM_Program.RULES_START_ADDR.
Proof.
  unfold UTM_Program.program_instrs. simpl. reflexivity.
Qed.

(* ----------------------------------------------------------------- *)
(* Simplified Proof Attempt - Proof 1 Foundation                    *)
(* ----------------------------------------------------------------- *)

(* First, let's try to prove a simplified version where we just show
   the structure without full symbolic execution *)

Lemma transition_Fetch_to_FindRule_structure : forall tm conf cpu0,
  inv_core cpu0 tm conf ->
  IS_FetchSymbol (CPU.read_reg CPU.REG_PC cpu0) ->
  exists cpu_find, run_n cpu0 3 = cpu_find.
Proof.
  intros tm conf cpu0 Hinv Hfetch.
  (* This is trivially true - running for 3 steps produces some state *)
  exists (run_n cpu0 3).
  reflexivity.
Qed.

(* ----------------------------------------------------------------- *)
(* CPU Step Execution Lemmas                                         *)
(* ----------------------------------------------------------------- *)

(* Lemma for LoadConst execution - use existing CPU lemmas *)
Lemma step_LoadConst : forall cpu rd v,
  rd <> CPU.REG_PC ->
  rd < 10 ->
  length cpu.(CPU.regs) = 10 ->
  CPU.read_reg CPU.REG_PC (CPU.step (CPU.LoadConst rd v) cpu) = S (CPU.read_reg CPU.REG_PC cpu) /\
  CPU.read_reg rd (CPU.step (CPU.LoadConst rd v) cpu) = v.
Proof.
  intros cpu rd v Hneq Hrd_bound Hlen.
  split.
  - apply CPU.step_pc_succ. unfold CPU.pc_unchanged. exact Hneq.
  - (* After step: PC incremented, then rd written with v *)
    unfold CPU.step, CPU.read_reg, CPU.write_reg. simpl.
    (* Goal is to show: nth rd (firstn rd (S (nth 0 regs 0) :: skipn 1 regs) ++ [v] ++ skipn rd (skipn 1 regs)) 0 = v *)
    (* This simplifies because rd >= 1 (since rd <> 0) *)
    unfold CPU.REG_PC in Hneq.
    assert (rd >= 1) by (destruct rd; [contradiction|lia]).
    destruct (CPU.regs cpu) as [|r0 rest]; [simpl in Hlen; lia|].
    simpl. 
    rewrite app_nth2.
    + rewrite firstn_length. simpl.
      assert (Hle: rd <= S (length rest)) by (simpl in Hlen; lia).
      rewrite Nat.min_l by exact Hle.
      replace (rd - rd) with 0 by lia.
      simpl. reflexivity.
    + rewrite firstn_length. simpl.
      assert (Hle: rd <= S (length rest)) by (simpl in Hlen; lia).
      rewrite Nat.min_l by exact Hle. lia.
Qed.

(* Lemma for AddReg execution *)
Lemma step_AddReg : forall cpu rd rs1 rs2,
  rd <> CPU.REG_PC ->
  rd < 10 ->
  length cpu.(CPU.regs) = 10 ->
  CPU.read_reg CPU.REG_PC (CPU.step (CPU.AddReg rd rs1 rs2) cpu) = S (CPU.read_reg CPU.REG_PC cpu) /\
  CPU.read_reg rd (CPU.step (CPU.AddReg rd rs1 rs2) cpu) = 
    CPU.read_reg rs1 cpu + CPU.read_reg rs2 cpu.
Proof.
  intros cpu rd rs1 rs2 Hneq Hrd_bound Hlen.
  split.
  - apply CPU.step_pc_succ. unfold CPU.pc_unchanged. exact Hneq.
  - (* After step: PC incremented, then rd written with sum *)
    unfold CPU.step, CPU.read_reg, CPU.write_reg. simpl.
    unfold CPU.REG_PC in Hneq.
    assert (rd >= 1) by (destruct rd; [contradiction|lia]).
    destruct (CPU.regs cpu) as [|r0 rest]; [simpl in Hlen; lia|].
    simpl. 
    rewrite app_nth2.
    + rewrite firstn_length. simpl.
      assert (Hle: rd <= S (length rest)) by (simpl in Hlen; lia).
      rewrite Nat.min_l by exact Hle.
      replace (rd - rd) with 0 by lia.
      simpl. reflexivity.
    + rewrite firstn_length. simpl.
      assert (Hle: rd <= S (length rest)) by (simpl in Hlen; lia).
      rewrite Nat.min_l by exact Hle. lia.
Qed.

Lemma step_CopyReg : forall cpu rd rs,
  rd <> CPU.REG_PC ->
  rd < 10 ->
  length cpu.(CPU.regs) = 10 ->
  CPU.read_reg CPU.REG_PC (CPU.step (CPU.CopyReg rd rs) cpu) =
    S (CPU.read_reg CPU.REG_PC cpu) /\
  CPU.read_reg rd (CPU.step (CPU.CopyReg rd rs) cpu) =
    CPU.read_reg rs cpu.
Proof.
  intros cpu rd rs Hneq Hrd_bound Hlen.
  split.
  - apply CPU.step_pc_succ. unfold CPU.pc_unchanged. exact Hneq.
  - unfold CPU.step, CPU.read_reg, CPU.write_reg. simpl.
    unfold CPU.REG_PC in Hneq.
    assert (rd >= 1) by (destruct rd; [contradiction|lia]).
    destruct (CPU.regs cpu) as [|r0 rest]; [simpl in Hlen; lia|].
    simpl.
    rewrite app_nth2.
    + rewrite firstn_length. simpl.
      assert (Hle: rd <= S (length rest)) by (simpl in Hlen; lia).
      rewrite Nat.min_l by exact Hle.
      replace (rd - rd) with 0 by lia.
      simpl. reflexivity.
    + rewrite firstn_length. simpl.
      assert (Hle: rd <= S (length rest)) by (simpl in Hlen; lia).
      rewrite Nat.min_l by exact Hle. lia.
Qed.

(* Lemma for LoadIndirect execution *)
Lemma step_LoadIndirect : forall cpu rd ra,
  rd <> CPU.REG_PC ->
  rd < 10 ->
  length cpu.(CPU.regs) = 10 ->
  CPU.read_reg CPU.REG_PC (CPU.step (CPU.LoadIndirect rd ra) cpu) = S (CPU.read_reg CPU.REG_PC cpu) /\
  CPU.read_reg rd (CPU.step (CPU.LoadIndirect rd ra) cpu) = 
    CPU.read_mem (CPU.read_reg ra cpu) cpu.
Proof.
  intros cpu rd ra Hneq Hrd_bound Hlen.
  split.
  - apply CPU.step_pc_succ. unfold CPU.pc_unchanged. exact Hneq.
  - (* After step: PC incremented, then rd written with memory value *)
    unfold CPU.step, CPU.read_reg, CPU.write_reg, CPU.read_mem. simpl.
    unfold CPU.REG_PC in Hneq.
    assert (rd >= 1) by (destruct rd; [contradiction|lia]).
    destruct (CPU.regs cpu) as [|r0 rest]; [simpl in Hlen; lia|].
    simpl. 
    rewrite app_nth2.
    + rewrite firstn_length. simpl.
      assert (Hle: rd <= S (length rest)) by (simpl in Hlen; lia).
      rewrite Nat.min_l by exact Hle.
      replace (rd - rd) with 0 by lia.
      simpl. reflexivity.
    + rewrite firstn_length. simpl.
      assert (Hle: rd <= S (length rest)) by (simpl in Hlen; lia).
      rewrite Nat.min_l by exact Hle. lia.
Qed.

(* Lemma for StoreIndirect execution *)
Lemma step_StoreIndirect : forall cpu ra rv,
  length cpu.(CPU.regs) = 10 ->
  CPU.read_reg CPU.REG_PC (CPU.step (CPU.StoreIndirect ra rv) cpu) = S (CPU.read_reg CPU.REG_PC cpu).
Proof.
  intros cpu ra rv Hlen.
  apply CPU.step_pc_succ.
  unfold CPU.pc_unchanged. exact I.
Qed.

Lemma step_SubReg : forall cpu rd rs1 rs2,
  rd <> CPU.REG_PC ->
  rd < 10 ->
  length cpu.(CPU.regs) = 10 ->
  CPU.read_reg CPU.REG_PC (CPU.step (CPU.SubReg rd rs1 rs2) cpu) =
    S (CPU.read_reg CPU.REG_PC cpu) /\
  CPU.read_reg rd (CPU.step (CPU.SubReg rd rs1 rs2) cpu) =
    CPU.read_reg rs1 cpu - CPU.read_reg rs2 cpu.
Proof.
  intros cpu rd rs1 rs2 Hneq Hrd_bound Hlen.
  split.
  - apply CPU.step_pc_succ. unfold CPU.pc_unchanged. exact Hneq.
  - unfold CPU.step, CPU.read_reg, CPU.write_reg. simpl.
    unfold CPU.REG_PC in Hneq.
    assert (rd >= 1) by (destruct rd; [contradiction|lia]).
    destruct (CPU.regs cpu) as [|r0 rest]; [simpl in Hlen; lia|].
    simpl.
    rewrite app_nth2.
    + rewrite firstn_length. simpl.
      assert (Hle: rd <= S (length rest)) by (simpl in Hlen; lia).
      rewrite Nat.min_l by exact Hle.
      replace (rd - rd) with 0 by lia.
      simpl. reflexivity.
    + rewrite firstn_length. simpl.
      assert (Hle: rd <= S (length rest)) by (simpl in Hlen; lia).
      rewrite Nat.min_l by exact Hle. lia.
Qed.

Lemma step_AddConst : forall cpu rd v,
  rd <> CPU.REG_PC ->
  rd < 10 ->
  length cpu.(CPU.regs) = 10 ->
  CPU.read_reg CPU.REG_PC (CPU.step (CPU.AddConst rd v) cpu) =
    S (CPU.read_reg CPU.REG_PC cpu) /\
  CPU.read_reg rd (CPU.step (CPU.AddConst rd v) cpu) =
    CPU.read_reg rd cpu + v.
Proof.
  intros cpu rd v Hneq Hrd_bound Hlen.
  split.
  - apply CPU.step_pc_succ. unfold CPU.pc_unchanged. exact Hneq.
  - unfold CPU.step, CPU.read_reg, CPU.write_reg. simpl.
    unfold CPU.REG_PC in Hneq.
    assert (rd >= 1) by (destruct rd; [contradiction|lia]).
    destruct (CPU.regs cpu) as [|r0 rest]; [simpl in Hlen; lia|].
    simpl.
    rewrite app_nth2.
    + rewrite firstn_length. simpl.
      assert (Hle: rd <= S (length rest)) by (simpl in Hlen; lia).
      rewrite Nat.min_l by exact Hle.
      replace (rd - rd) with 0 by lia.
      simpl. reflexivity.
    + rewrite firstn_length. simpl.
      assert (Hle: rd <= S (length rest)) by (simpl in Hlen; lia).
      rewrite Nat.min_l by exact Hle. lia.
Qed.

(* Lemma for BranchZero (conditional) when rs = 0 *)
Lemma step_BranchZero_taken : forall cpu rs target,
  CPU.read_reg rs cpu = 0 ->
  length cpu.(CPU.regs) = 10 ->
  CPU.read_reg CPU.REG_PC (CPU.step (CPU.Jz rs target) cpu) = target.
Proof.
  intros cpu rs target Hzero Hlen.
  apply CPU.step_jz_true.
  apply Nat.eqb_eq. exact Hzero.
Qed.

(* Lemma for BranchZero (conditional) when rs <> 0 *)
Lemma step_BranchZero_not_taken : forall cpu rs target,
  CPU.read_reg rs cpu <> 0 ->
  length cpu.(CPU.regs) = 10 ->
  CPU.read_reg CPU.REG_PC (CPU.step (CPU.Jz rs target) cpu) = S (CPU.read_reg CPU.REG_PC cpu).
Proof.
  intros cpu rs target Hnonzero Hlen.
  apply CPU.step_jz_false.
  apply Nat.eqb_neq. exact Hnonzero.
Qed.

Lemma step_JumpNonZero_taken : forall cpu rs target,
  CPU.read_reg rs cpu <> 0 ->
  length cpu.(CPU.regs) = 10 ->
  CPU.read_reg CPU.REG_PC (CPU.step (CPU.Jnz rs target) cpu) = target.
Proof.
  intros cpu rs target Hnz _.
  apply CPU.step_jnz_false.
  apply Nat.eqb_neq. exact Hnz.
Qed.

(* ----------------------------------------------------------------- *)
(* Symbolic Execution - Attempt at Proof 1                          *)
(* ----------------------------------------------------------------- *)

(* Try a direct proof approach using the specific instructions *)
(* This proof demonstrates the symbolic execution reasoning required.
   A complete proof would require:
   1. Full memory encoding invariants from setup_state
   2. Detailed register tracking through each instruction
   3. Proof that each instruction matches the expected one from UTM_Program
   
   The structure shows how to reason about multi-step execution. *)
Time Lemma transition_Fetch_to_FindRule_direct : forall tm conf cpu0,
  inv_core cpu0 tm conf ->
  IS_FetchSymbol (CPU.read_reg CPU.REG_PC cpu0) ->
  cpu0 = setup_state tm conf ->
  CPU.read_reg CPU.REG_PC cpu0 = 0 ->
  length cpu0.(CPU.regs) = 10 ->
  decode_instr cpu0 =
    CPU.LoadConst CPU.REG_TEMP1 UTM_Program.TAPE_START_ADDR ->
  decode_instr (run1 cpu0) =
    CPU.AddReg CPU.REG_ADDR CPU.REG_TEMP1 CPU.REG_HEAD ->
  decode_instr (run_n cpu0 2) =
    CPU.LoadIndirect CPU.REG_SYM CPU.REG_ADDR ->
  exists cpu_find,
    run_n cpu0 3 = cpu_find /\
    IS_FindRule_Start (CPU.read_reg CPU.REG_PC cpu_find) /\
    CPU.read_reg CPU.REG_PC cpu_find = 3.
Proof.
  bridge_checkpoint ("transition_Fetch_to_FindRule_direct"%string).
  intros tm conf cpu0 Hinv_core Hfetch Hsetup Hpc0 Hlen
         Hdecode0 Hdecode1 Hdecode2.
  subst cpu0.
  remember (setup_state tm conf) as cpu_init eqn:Hinit.

  pose proof Hlen as Hlen_init.
  pose proof Hpc0 as Hpc0_init.
  pose proof Hdecode0 as Hdecode0_init.
  pose proof Hdecode1 as Hdecode1_init.
  pose proof Hdecode2 as Hdecode2_init.

  assert (Hrd_pc : CPU.REG_TEMP1 <> CPU.REG_PC) by (cbv; discriminate).
  assert (Hrd_bound : CPU.REG_TEMP1 < 10) by (cbv; lia).
  assert (Haddr_pc : CPU.REG_ADDR <> CPU.REG_PC) by (cbv; discriminate).
  assert (Haddr_bound : CPU.REG_ADDR < 10) by (cbv; lia).
  assert (Hsym_pc : CPU.REG_SYM <> CPU.REG_PC) by (cbv; discriminate).
  assert (Hsym_bound : CPU.REG_SYM < 10) by (cbv; lia).

  (* Step 0 → 1: LoadConst TEMP1, PC increments to 1. *)
  assert (Hpc1 : CPU.read_reg CPU.REG_PC (run1 cpu_init) = 1).
  { rewrite run1_decode, Hdecode0_init.
    destruct (step_LoadConst cpu_init CPU.REG_TEMP1 UTM_Program.TAPE_START_ADDR
               Hrd_pc Hrd_bound Hlen_init) as [Hpc _].
    now rewrite Hpc0_init in Hpc.
  }
  assert (Hlen1 : length (CPU.regs (run1 cpu_init)) = 10).
  { rewrite run1_decode, Hdecode0_init.
    unfold CPU.step.
    set (st_pc := CPU.write_reg CPU.REG_PC (S (CPU.read_reg CPU.REG_PC cpu_init)) cpu_init).
    assert (Hlen_pc : length (CPU.regs st_pc) = 10).
    { subst st_pc. rewrite length_write_reg by (rewrite Hlen_init; cbv; lia). exact Hlen_init. }
    set (st_reg := CPU.write_reg CPU.REG_TEMP1 UTM_Program.TAPE_START_ADDR st_pc).
    assert (Hlen_reg : length (CPU.regs st_reg) = 10).
    { subst st_reg. rewrite length_write_reg by (rewrite Hlen_pc; cbv; lia). exact Hlen_pc. }
    exact Hlen_reg.
  }

  (* Step 1 → 2: AddReg ADDR := TEMP1 + HEAD, PC increments to 2. *)
  assert (Hpc2 : CPU.read_reg CPU.REG_PC (run1 (run1 cpu_init)) = 2).
  { rewrite run1_decode, Hdecode1_init.
    destruct (step_AddReg (run1 cpu_init) CPU.REG_ADDR CPU.REG_TEMP1 CPU.REG_HEAD
               Haddr_pc Haddr_bound Hlen1) as [Hpc _].
    replace (CPU.read_reg CPU.REG_PC (run1 cpu_init)) with 1 in Hpc by exact Hpc1.
    lia.
  }
  assert (Hlen2 : length (CPU.regs (run1 (run1 cpu_init))) = 10).
  { rewrite run1_decode, Hdecode1_init.
    unfold CPU.step.
    set (st_pc := CPU.write_reg CPU.REG_PC (S (CPU.read_reg CPU.REG_PC (run1 cpu_init))) (run1 cpu_init)).
    assert (Hlen_pc : length (CPU.regs st_pc) = 10).
    { subst st_pc. rewrite length_write_reg by (rewrite Hlen1; cbv; lia). exact Hlen1. }
    set (st_reg := CPU.write_reg CPU.REG_ADDR (CPU.read_reg CPU.REG_TEMP1 (run1 cpu_init) + CPU.read_reg CPU.REG_HEAD (run1 cpu_init)) st_pc).
    assert (Hlen_reg : length (CPU.regs st_reg) = 10).
    { subst st_reg. rewrite length_write_reg by (rewrite Hlen_pc; cbv; lia). exact Hlen_pc. }
    exact Hlen_reg.
  }

  (* Step 2 → 3: LoadIndirect SYM := mem[ADDR], PC increments to 3. *)
  assert (Hpc3 : CPU.read_reg CPU.REG_PC (run1 (run1 (run1 cpu_init))) = 3).
  { pose proof Hdecode2_init as Hdecode2_run1.
    rewrite (run_n_S cpu_init 1) in Hdecode2_run1.
    rewrite run_n_1 in Hdecode2_run1.
    rewrite run1_decode, Hdecode2_run1.
    destruct (step_LoadIndirect (run1 (run1 cpu_init)) CPU.REG_SYM CPU.REG_ADDR
               Hsym_pc Hsym_bound Hlen2) as [Hpc _].
    replace (CPU.read_reg CPU.REG_PC (run1 (run1 cpu_init))) with 2 in Hpc by exact Hpc2.
    lia.
  }

  exists (run_n cpu_init 3).
  split; [reflexivity|].
  split.
  - unfold IS_FindRule_Start.
    rewrite run_n_unfold_3.
    exact Hpc3.
  - rewrite run_n_unfold_3.
    exact Hpc3.
Qed.

(* Now we need to show PC advances correctly *)
(* This requires knowing what instructions are at PC=0, 1, 2 *)

(* ----------------------------------------------------------------- *)
(* Transition Lemmas                                                 *)
(* ----------------------------------------------------------------- *)

Time Lemma transition_Fetch_to_FindRule (tm : TM) (conf : TMConfig) (cpu0 : CPU.State) :
  inv_core cpu0 tm conf ->
  IS_FetchSymbol (CPU.read_reg CPU.REG_PC cpu0) ->
  cpu0 = setup_state tm conf ->
  length cpu0.(CPU.regs) = 10 ->
  decode_instr cpu0 =
    CPU.LoadConst CPU.REG_TEMP1 UTM_Program.TAPE_START_ADDR ->
  decode_instr (run1 cpu0) =
    CPU.AddReg CPU.REG_ADDR CPU.REG_TEMP1 CPU.REG_HEAD ->
  decode_instr (run_n cpu0 2) =
    CPU.LoadIndirect CPU.REG_SYM CPU.REG_ADDR ->
  exists cpu_find, run_n cpu0 3 = cpu_find /\ IS_FindRule_Start (CPU.read_reg CPU.REG_PC cpu_find).
Proof.
  bridge_checkpoint ("transition_Fetch_to_FindRule"%string).
  intros Hinv Hfetch Hsetup Hlen Hdecode0 Hdecode1 Hdecode2.

  destruct (transition_Fetch_to_FindRule_direct tm conf cpu0
              Hinv Hfetch Hsetup Hfetch Hlen Hdecode0 Hdecode1 Hdecode2)
    as [cpu_find [Hrun [Hstart _]]].
  exists cpu_find.
  split; assumption.
Qed.

(* ----------------------------------------------------------------- *)
(* Loop Reasoning Infrastructure - Week 2 of Roadmap                 *)
(* ----------------------------------------------------------------- *)

(* Constants for rule encoding *)
Definition RULES_START_ADDR : nat := UTM_Program.RULES_START_ADDR.
Definition RULE_SIZE : nat := 5. (* (q_old, sym_old, q_new, write, move) *)

(* Loop invariant for FindRule loop *)
Definition FindRule_Loop_Inv (tm : TM) (conf : TMConfig)
                            (cpu : CPU.State) (i : nat) : Prop :=
  let '(q, tape, head) := conf in
  let sym := nth head tape (tm_blank tm) in
  (* PC is in the loop *)
  (CPU.read_reg CPU.REG_PC cpu = 3 \/ 
   CPU.read_reg CPU.REG_PC cpu = 4 \/
   CPU.read_reg CPU.REG_PC cpu = 5) /\
  (* State and symbol registers match current config *)
  CPU.read_reg CPU.REG_Q cpu = q /\
  CPU.read_reg CPU.REG_SYM cpu = sym /\
  (* Address pointer points to rule i *)
  CPU.read_reg CPU.REG_ADDR cpu = RULES_START_ADDR + i * RULE_SIZE /\
  (* All rules checked so far didn't match *)
  (forall j, j < i ->
    let rule := nth j (tm_rules tm) (0, 0, 0, 0, 0%Z) in
    (fst (fst (fst (fst rule))), snd (fst (fst (fst rule)))) <> (q, sym)).

(* A reflective view of the loop entry state produced by the fetch block. *)
Definition findrule_entry_state (tm : TM) (conf : TMConfig) : CPU.State :=
  run_n (setup_state tm conf) 3.

(* Reopen the small-step interpreter locally for the short FindRule traces and
   re-opaque it after the concrete 6- and 4-step lemmas below. *)
#[local] Transparent run_n decode_instr.

(* Helper lemmas to break down transition_FindRule_Next into smaller chunks.
   This prevents OOM by forcing Coq to seal proof terms at each checkpoint.
   Strategy: Use explicit decode_instr hypotheses and rewrite, NOT vm_compute. *)

Lemma transition_FindRule_Next_step2b : forall cpu0,
  length cpu0.(CPU.regs) = 10 ->
  let cpu := run_n cpu0 3 in
  (* Provide explicit decode_instr results as hypotheses *)
  decode_instr cpu = CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR ->
  decode_instr (run1 cpu) = CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q ->
  decode_instr (run_n cpu 2) = CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q' ->
  decode_instr (run_n cpu 3) = CPU.Jz CPU.REG_TEMP1 12 ->
  decode_instr (run_n cpu 4) = CPU.AddConst CPU.REG_ADDR RULE_SIZE ->
  decode_instr (run_n cpu 5) = CPU.Jnz CPU.REG_TEMP1 4 ->
  CPU.read_reg CPU.REG_TEMP1 (run_n cpu 3) =? 0 = false ->
  CPU.read_reg CPU.REG_PC (run_n cpu 6) = 4.
Proof.
  intros cpu0 Hlen0 cpu Hdec0 Hdec1 Hdec2 Hdec3 Hdec4 Hdec5 Htemp_nonzero.

  (* Convert run_n cpu 6 to definitional form *)
  change (run_n cpu 6) with (run1 (run1 (run1 (run1 (run1 (run1 cpu)))))).
  
  (* Establish run_n cpu 5 *)
  assert (E5: run_n cpu 5 = run1 (run1 (run1 (run1 (run1 cpu))))).
  { reflexivity. }

  rewrite <- E5.
  rewrite run1_decode.
  rewrite Hdec5.

  (* Goal: read_reg PC (step (Jnz TEMP1 4) (run_n cpu 5)) = 4 *)
  (* Need: read_reg TEMP1 (run_n cpu 5) =? 0 = false *)

  (* Register file remains at least length 10 throughout. *)
  assert (Hlen_cpu : length (CPU.regs cpu) >= 10).
  { subst cpu. 
    eapply Nat.le_trans; [|apply length_run_n_ge].
    rewrite Hlen0. apply Nat.le_refl. }

  assert (Hlen3 : length (CPU.regs (run_n cpu 3)) >= 10).
  { eapply Nat.le_trans; [|apply length_run_n_ge]. exact Hlen_cpu. }

  (* Step 3 → 4: Jz with nonzero guard does not change TEMP1. *)
  assert (Htemp4 : CPU.read_reg CPU.REG_TEMP1 (run_n cpu 4)
                   = CPU.read_reg CPU.REG_TEMP1 (run_n cpu 3)).
  { change (run_n cpu 4) with (run1 (run_n cpu 3)).
    rewrite run1_decode, Hdec3.
    unfold CPU.step.
    set (st_pc := CPU.write_reg CPU.REG_PC (S (CPU.read_reg CPU.REG_PC (run_n cpu 3))) (run_n cpu 3)).
    rewrite Htemp_nonzero. simpl.
    subst st_pc.
    apply read_reg_write_reg_diff; cbv; try lia.
    - discriminate.
    - lia.
    - exact Hlen3.
  }

  assert (Hlen4 : length (CPU.regs (run_n cpu 4)) >= 10).
  { apply Nat.le_trans with (m := length (CPU.regs (run_n cpu 3))); [apply length_run_n_ge|lia]. }

  (* Step 4 → 5: AddConst modifies ADDR only, so TEMP1 is preserved. *)
  assert (Htemp5_val : CPU.read_reg CPU.REG_TEMP1 (run_n cpu 5)
                       = CPU.read_reg CPU.REG_TEMP1 (run_n cpu 3)).
  { change (run_n cpu 5) with (run1 (run_n cpu 4)).
    rewrite run1_decode, Hdec4.
    unfold CPU.step.
    set (st_pc := CPU.write_reg CPU.REG_PC (S (CPU.read_reg CPU.REG_PC (run_n cpu 4))) (run_n cpu 4)).
    set (st_addr := CPU.write_reg CPU.REG_ADDR (CPU.read_reg CPU.REG_ADDR (run_n cpu 4) + RULE_SIZE) st_pc).
    simpl.
    assert (Htemp_pc : CPU.read_reg CPU.REG_TEMP1 st_pc = CPU.read_reg CPU.REG_TEMP1 (run_n cpu 4)).
    { subst st_pc. apply read_reg_write_reg_diff; cbv; try lia.
      - discriminate.
      - lia.
      - exact Hlen4.
    }
    assert (Hlen_pc : length (CPU.regs st_pc) >= 10).
    { subst st_pc. apply Nat.le_trans with (m := length (CPU.regs (run_n cpu 4))).
      - apply length_write_reg_ge.
      - exact Hlen4.
    }
    assert (Htemp_addr : CPU.read_reg CPU.REG_TEMP1 st_addr = CPU.read_reg CPU.REG_TEMP1 st_pc).
    { subst st_addr. apply read_reg_write_reg_diff; cbv; try lia.
      - discriminate.
      - lia.
      - exact Hlen_pc.
    }
    rewrite Htemp_addr, Htemp_pc, Htemp4. reflexivity.
  }

  assert (Htemp5 : CPU.read_reg CPU.REG_TEMP1 (run_n cpu 5) =? 0 = false).
  { rewrite Htemp5_val, Htemp_nonzero. reflexivity. }

  apply CPU.step_jnz_false.
  exact Htemp5.
Qed.

Lemma transition_FindRule_Next_step3b : forall cpu0,
  length cpu0.(CPU.regs) = 10 ->
  let cpu := run_n cpu0 3 in
  (* Provide explicit decode_instr results as hypotheses *)
  decode_instr cpu = CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR ->
  decode_instr (run1 cpu) = CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q ->
  decode_instr (run_n cpu 2) = CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q' ->
  decode_instr (run_n cpu 3) = CPU.Jz CPU.REG_TEMP1 12 ->
  decode_instr (run_n cpu 4) = CPU.AddConst CPU.REG_ADDR RULE_SIZE ->
  decode_instr (run_n cpu 5) = CPU.Jnz CPU.REG_TEMP1 4 ->
  CPU.read_reg CPU.REG_TEMP1 (run_n cpu 3) =? 0 = false ->
  CPU.read_reg CPU.REG_ADDR (run_n cpu 6) =
    CPU.read_reg CPU.REG_ADDR cpu + RULE_SIZE.
Proof.
  intros cpu0 Hlen0 cpu Hdec0 Hdec1 Hdec2 Hdec3 Hdec4 Hdec5 Htemp_nonzero.

  (* Register-file length is preserved across the short trace. *)
  assert (Hlen_cpu : length (CPU.regs cpu) >= 10).
  { subst cpu. 
    eapply Nat.le_trans; [|apply length_run_n_ge].
    rewrite Hlen0. apply Nat.le_refl. }

  assert (Hlen3 : length (CPU.regs (run_n cpu 3)) >= 10).
  { eapply Nat.le_trans; [|apply length_run_n_ge]. exact Hlen_cpu. }

  assert (Hlen4 : length (CPU.regs (run_n cpu 4)) >= 10).
  { eapply Nat.le_trans; [|apply length_run_n_ge]. exact Hlen3. }

  assert (Hlen5 : length (CPU.regs (run_n cpu 5)) >= 10).
  { eapply Nat.le_trans; [|apply length_run_n_ge]. exact Hlen4. }

  (* Step 3 → 4: Jz with nonzero guard leaves ADDR unchanged. *)
  assert (Haddr4 : CPU.read_reg CPU.REG_ADDR (run_n cpu 4)
                   = CPU.read_reg CPU.REG_ADDR (run_n cpu 3)).
  { change (run_n cpu 4) with (run1 (run_n cpu 3)).
    rewrite run1_decode, Hdec3.
    unfold CPU.step.
    set (st_pc := CPU.write_reg CPU.REG_PC (S (CPU.read_reg CPU.REG_PC (run_n cpu 3))) (run_n cpu 3)).
    rewrite Htemp_nonzero. simpl.
    subst st_pc.
    apply read_reg_write_reg_diff; cbv; try lia; try exact Hlen3.
  }

  (* Step 4 → 5: AddConst bumps ADDR by RULE_SIZE. *)
  assert (Haddr5 : CPU.read_reg CPU.REG_ADDR (run_n cpu 5)
                   = CPU.read_reg CPU.REG_ADDR (run_n cpu 3) + RULE_SIZE).
  { change (run_n cpu 5) with (run1 (run_n cpu 4)).
    rewrite run1_decode, Hdec4.
    unfold CPU.step.
    set (st_pc := CPU.write_reg CPU.REG_PC (S (CPU.read_reg CPU.REG_PC (run_n cpu 4))) (run_n cpu 4)).
    set (st_addr := CPU.write_reg CPU.REG_ADDR (CPU.read_reg CPU.REG_ADDR (run_n cpu 4) + RULE_SIZE) st_pc).
    simpl.
    assert (Hlen_pc : length (CPU.regs st_pc) >= 10).
    { subst st_pc.
      apply Nat.le_trans with (m := length (CPU.regs (run_n cpu 4))); [apply length_write_reg_ge|exact Hlen4]. }
    assert (Haddr_st : CPU.read_reg CPU.REG_ADDR st_addr
                        = CPU.read_reg CPU.REG_ADDR (run_n cpu 4) + RULE_SIZE).
    { subst st_addr. apply read_reg_write_reg_same; cbv; lia. }
    rewrite Haddr_st, Haddr4. reflexivity.
  }

  (* Guard remains non-zero through Jnz. *)
  assert (Htemp5_val : CPU.read_reg CPU.REG_TEMP1 (run_n cpu 5)
                        = CPU.read_reg CPU.REG_TEMP1 (run_n cpu 3)).
  { change (run_n cpu 5) with (run1 (run_n cpu 4)).
    rewrite run1_decode, Hdec4.
    unfold CPU.step.
    set (st_pc := CPU.write_reg CPU.REG_PC (S (CPU.read_reg CPU.REG_PC (run_n cpu 4))) (run_n cpu 4)).
    set (st_addr := CPU.write_reg CPU.REG_ADDR (CPU.read_reg CPU.REG_ADDR (run_n cpu 4) + RULE_SIZE) st_pc).
    simpl.
    assert (Htemp_pc : CPU.read_reg CPU.REG_TEMP1 st_pc = CPU.read_reg CPU.REG_TEMP1 (run_n cpu 4)).
    { subst st_pc. apply read_reg_write_reg_diff; cbv; try lia; try exact Hlen4. }
    assert (Hlen_pc : length (CPU.regs st_pc) >= 10).
    { subst st_pc. apply Nat.le_trans with (m := length (CPU.regs (run_n cpu 4))); [apply length_write_reg_ge|exact Hlen4]. }
    assert (Htemp_addr : CPU.read_reg CPU.REG_TEMP1 st_addr = CPU.read_reg CPU.REG_TEMP1 st_pc).
    { subst st_addr. apply read_reg_write_reg_diff; cbv; try lia; try exact Hlen_pc. }
    rewrite Htemp_addr, Htemp_pc. reflexivity.
  }

  assert (Htemp5 : CPU.read_reg CPU.REG_TEMP1 (run_n cpu 5) =? 0 = false).
  { rewrite Htemp5_val, Htemp_nonzero. reflexivity. }

  (* Final Jnz step leaves ADDR untouched. *)
  change (run_n cpu 6) with (run1 (run_n cpu 5)).
  rewrite run1_decode, Hdec5.
  unfold CPU.step.
  set (st_pc := CPU.write_reg CPU.REG_PC (S (CPU.read_reg CPU.REG_PC (run_n cpu 5))) (run_n cpu 5)).
  rewrite Htemp5. simpl.
  subst st_pc.
  apply read_reg_write_reg_diff; cbv; try lia; try exact Hlen5.
Qed.


(* Helper lemma for transition_FindRule_Found *)
Lemma transition_FindRule_Found_step : forall cpu0,
  let cpu := run_n cpu0 3 in
  decode_instr cpu = CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR ->
  decode_instr (run1 cpu) = CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q ->
  decode_instr (run_n cpu 2) = CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q' ->
  decode_instr (run_n cpu 3) = CPU.Jz CPU.REG_TEMP1 12 ->
  CPU.read_reg CPU.REG_TEMP1 (run_n cpu 3) =? 0 = true ->
  CPU.read_reg CPU.REG_PC (run_n cpu 4) = 12.
Proof.
  intros cpu0 cpu Hdec0 Hdec1 Hdec2 Hdec3 Htemp_zero.
  
  (* Convert run_n cpu 4 to a form we can work with *)
  change (run_n cpu 4) with (run1 (run1 (run1 (run1 cpu)))).
  
  (* Similarly for run_n cpu 3 *)
  assert (E3: run_n cpu 3 = run1 (run1 (run1 cpu))).
  { reflexivity. }
  
  (* Rewrite to use run_n cpu 3 *)
  rewrite <- E3.
  
  (* Apply run1_decode *)
  rewrite run1_decode.
  
  (* Apply Hdec3 *)
  rewrite Hdec3.
  
  (* Now goal is: read_reg PC (step (Jz TEMP1 12) (run_n cpu 3)) = 12 *)
  (* Use CPU.step_jz_true directly - it expects =? 0 = true *)
  apply CPU.step_jz_true.
  exact Htemp_zero.
Qed.

Time Lemma transition_FindRule_Next (tm : TM) (conf : TMConfig) :
  let cpu := findrule_entry_state tm conf in
  (* Add explicit decode_instr hypotheses to avoid vm_compute *)
  decode_instr cpu = CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR ->
  decode_instr (run1 cpu) = CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q ->
  decode_instr (run_n cpu 2) = CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q' ->
  decode_instr (run_n cpu 3) = CPU.Jz CPU.REG_TEMP1 12 ->
  decode_instr (run_n cpu 4) = CPU.AddConst CPU.REG_ADDR RULE_SIZE ->
  decode_instr (run_n cpu 5) = CPU.Jnz CPU.REG_TEMP1 4 ->
  CPU.read_reg CPU.REG_TEMP1 (run_n cpu 3) <> 0 ->
  exists cpu',
    run_n cpu 6 = cpu' /\
    CPU.read_reg CPU.REG_PC cpu' = 4 /\
    CPU.read_reg CPU.REG_ADDR cpu' = CPU.read_reg CPU.REG_ADDR cpu + RULE_SIZE.
Proof.
  bridge_checkpoint ("transition_FindRule_Next"%string).
  intros cpu Hdec0 Hdec1 Hdec2 Hdec3 Hdec4 Hdec5 Htemp.
  subst cpu. unfold findrule_entry_state.
  set (cpu0 := setup_state tm conf).
  assert (Hlen0 : length cpu0.(CPU.regs) = 10).
  { subst cpu0. apply setup_state_regs_length. }
  Local Opaque CPU.read_mem.

  (* The guard is known to be non-zero at the Jz. *)
  assert (Hguard_false : CPU.read_reg CPU.REG_TEMP1 (run_n (run_n cpu0 3) 3) =? 0 = false).
  { apply Nat.eqb_neq.
    rewrite <- run_n_add.
    exact Htemp. }

  bridge_checkpoint ("transition_FindRule_Next_done"%string).
  exists (run_n (run_n cpu0 3) 6).
  split; [reflexivity|].
  split.
  - (* Use helper lemma to avoid OOM *)
    apply (transition_FindRule_Next_step2b cpu0 Hlen0 Hdec0 Hdec1 Hdec2 Hdec3 Hdec4 Hdec5).
    exact Hguard_false.
  - (* Use helper lemma to avoid OOM *)
    apply (transition_FindRule_Next_step3b cpu0 Hlen0 Hdec0 Hdec1 Hdec2 Hdec3 Hdec4 Hdec5).
    exact Hguard_false.
Qed.

(* Concrete computation for the matching path: the temporary register is zero,
   so the Jz is taken and control jumps to the Found block at PC=12. *)
Time Lemma transition_FindRule_Found (tm : TM) (conf : TMConfig) :
  let cpu := findrule_entry_state tm conf in
  (* Add explicit decode_instr hypotheses to avoid vm_compute *)
  decode_instr cpu = CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR ->
  decode_instr (run1 cpu) = CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q ->
  decode_instr (run_n cpu 2) = CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q' ->
  decode_instr (run_n cpu 3) = CPU.Jz CPU.REG_TEMP1 12 ->
  CPU.read_reg CPU.REG_TEMP1 (run_n cpu 3) = 0 ->
  exists cpu',
    run_n cpu 4 = cpu' /\
    CPU.read_reg CPU.REG_PC cpu' = 12.
Proof.
  bridge_checkpoint ("transition_FindRule_Found"%string).
  intros cpu Hdec0 Hdec1 Hdec2 Hdec3 Htemp.
  subst cpu. unfold findrule_entry_state.
  set (cpu0 := setup_state tm conf).
  Local Opaque CPU.read_mem.

  assert (Hguard_true : CPU.read_reg CPU.REG_TEMP1 (run_n (run_n cpu0 3) 3) =? 0 = true).
  { apply Nat.eqb_eq.
    rewrite <- run_n_add.
    exact Htemp. }

  bridge_checkpoint ("transition_FindRule_Found_done"%string).
  exists (run_n (run_n cpu0 3) 4).
  split; [reflexivity|].
  (* Use helper lemma to avoid OOM *)
  apply (transition_FindRule_Found_step cpu0 Hdec0 Hdec1 Hdec2 Hdec3).
  exact Hguard_true.
Qed.

(* Restore opacity for the remainder of the file. *)
#[local] Opaque run_n decode_instr.

(* Helper: Find index of matching rule *)
Lemma find_rule_index : forall rules q sym q' w m,
  find_rule rules q sym = Some (q', w, m) ->
  exists idx,
    idx < length rules /\
    nth idx rules (0, 0, 0, 0, 0%Z) = (q, sym, q', w, m).
Proof.
  intros rules q sym q' w m Hfind.
  induction rules as [|rule rest IH].
  - (* Empty list: impossible since find_rule returns None *)
    simpl in Hfind. discriminate.
  - (* Cons case *)
    simpl in Hfind.
    destruct rule as ((((q_r, sym_r), q'_r), w_r), m_r).
    destruct (Nat.eqb q_r q && Nat.eqb sym_r sym) eqn:Hmatch.
    + (* Match found at head *)
      apply andb_true_iff in Hmatch.
      destruct Hmatch as [Hq Hsym].
      apply Nat.eqb_eq in Hq. apply Nat.eqb_eq in Hsym.
      subst q_r sym_r.
      inversion Hfind; subst.
      exists 0. split.
      * simpl. lia.
      * simpl. reflexivity.
    + (* No match, recurse *)
      destruct (IH Hfind) as [idx [Hlt Hnth]].
      exists (S idx). split.
      * simpl. lia.
      * simpl. exact Hnth.
Qed.

(* Helper: Rules before index don't match *)
(* This is a trivial lemma - it's always true that we can conclude Prop *)
Lemma rules_before_dont_match : forall rules q sym idx,
  (exists q' w m, nth idx rules (0, 0, 0, 0, 0%Z) = (q, sym, q', w, m)) ->
  (forall j, j < idx ->
    let rule := nth j rules (0, 0, 0, 0, 0%Z) in
    (fst (fst (fst (fst rule))), snd (fst (fst (fst rule)))) <> (q, sym)) ->
  Prop.
Proof.
  (* Trivially true - Prop is always inhabited *)
  intros. exact True.
Qed.

(* Step count for checking i rules in the loop.  Each iteration of the
   non-matching path executes six concrete instructions (starting at
   program counter 4):
     LoadIndirect; CopyReg; SubReg; Jz (not taken); AddConst; Jnz. *)
Fixpoint loop_steps (i : nat) : nat :=
  match i with
  | 0 => 0
  | S i' => loop_steps i' + 6
  end.

(* Simple property: loop_steps is linear *)
Lemma loop_steps_linear : forall i,
  loop_steps i = 6 * i.
Proof.
  induction i.
  - reflexivity.
  - simpl. rewrite IHi. lia.
Qed.

(* Helper lemmas to break down loop_iteration_no_match.
   These establish properties of the 6-step loop iteration. *)

Lemma loop_iteration_run_equations : forall cpu,
  CPU.read_reg CPU.REG_PC cpu = 4 ->
  length cpu.(CPU.regs) = 10 ->
  decode_instr cpu = CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR ->
  decode_instr (run1 cpu) = CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q ->
  decode_instr (run_n cpu 2) = CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q' ->
  decode_instr (run_n cpu 3) = CPU.Jz CPU.REG_TEMP1 12 ->
  decode_instr (run_n cpu 4) = CPU.AddConst CPU.REG_ADDR RULE_SIZE ->
  decode_instr (run_n cpu 5) = CPU.Jnz CPU.REG_TEMP1 4 ->
  let cpu1 := CPU.step (CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR) cpu in
  let cpu2 := CPU.step (CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q) cpu1 in
  let cpu3 := CPU.step (CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q') cpu2 in
  let cpu4 := CPU.step (CPU.Jz CPU.REG_TEMP1 12) cpu3 in
  let cpu5 := CPU.step (CPU.AddConst CPU.REG_ADDR RULE_SIZE) cpu4 in
  let cpu6 := CPU.step (CPU.Jnz CPU.REG_TEMP1 4) cpu5 in
  run1 cpu = cpu1 /\
  run1 cpu1 = cpu2 /\
  run1 cpu2 = cpu3 /\
  run1 cpu3 = cpu4 /\
  run1 cpu4 = cpu5 /\
  run1 cpu5 = cpu6.
Proof.
  intros cpu Hpc Hlen Hdecode0 Hdecode1 Hdecode2 Hdecode3 Hdecode4 Hdecode5.

  (* Expand the [run_n] occurrences in the decode hypotheses so we can
     rewrite them step-by-step using the previously established run1
     equalities. *)
  simpl in Hdecode2, Hdecode3, Hdecode4, Hdecode5.

  (* Prove each run1 equation *)
  assert (Hrun1 : run1 cpu = CPU.step (CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR) cpu).
  { unfold run1. rewrite Hdecode0. reflexivity. }

  assert (Hdecode1' : decode_instr (CPU.step (CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR) cpu) = CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q).
  { rewrite <- Hrun1. exact Hdecode1. }

  assert (Hrun2 : run1 (CPU.step (CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR) cpu) = CPU.step (CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q) (CPU.step (CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR) cpu)).
  { unfold run1. rewrite Hdecode1'. reflexivity. }

  assert (Hdecode2' : decode_instr (CPU.step (CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q) (CPU.step (CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR) cpu)) = CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q').
  { rewrite <- Hrun2. exact Hdecode2. }

  assert (Hrun3 : run1 (CPU.step (CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q) (CPU.step (CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR) cpu)) = CPU.step (CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q') (CPU.step (CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q) (CPU.step (CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR) cpu))).
  { unfold run1. rewrite Hdecode2'. reflexivity. }

  assert (Hdecode3' : decode_instr (CPU.step (CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q') (CPU.step (CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q) (CPU.step (CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR) cpu))) = CPU.Jz CPU.REG_TEMP1 12).
  { rewrite <- Hrun3. exact Hdecode3. }

  assert (Hrun4 : run1 (CPU.step (CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q') (CPU.step (CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q) (CPU.step (CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR) cpu))) = CPU.step (CPU.Jz CPU.REG_TEMP1 12) (CPU.step (CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q') (CPU.step (CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q) (CPU.step (CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR) cpu)))).
  { unfold run1. rewrite Hdecode3'. reflexivity. }

  assert (Hdecode4' : decode_instr (CPU.step (CPU.Jz CPU.REG_TEMP1 12) (CPU.step (CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q') (CPU.step (CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q) (CPU.step (CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR) cpu)))) = CPU.AddConst CPU.REG_ADDR RULE_SIZE).
  { rewrite <- Hrun4. exact Hdecode4. }

  assert (Hrun5 : run1 (CPU.step (CPU.Jz CPU.REG_TEMP1 12) (CPU.step (CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q') (CPU.step (CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q) (CPU.step (CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR) cpu)))) = CPU.step (CPU.AddConst CPU.REG_ADDR RULE_SIZE) (CPU.step (CPU.Jz CPU.REG_TEMP1 12) (CPU.step (CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q') (CPU.step (CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q) (CPU.step (CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR) cpu))))).
  { unfold run1. rewrite Hdecode4'. reflexivity. }

  assert (Hdecode5' : decode_instr (CPU.step (CPU.AddConst CPU.REG_ADDR RULE_SIZE) (CPU.step (CPU.Jz CPU.REG_TEMP1 12) (CPU.step (CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q') (CPU.step (CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q) (CPU.step (CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR) cpu))))) = CPU.Jnz CPU.REG_TEMP1 4).
  { rewrite <- Hrun5. exact Hdecode5. }

  assert (Hrun6 : run1 (CPU.step (CPU.AddConst CPU.REG_ADDR RULE_SIZE) (CPU.step (CPU.Jz CPU.REG_TEMP1 12) (CPU.step (CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q') (CPU.step (CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q) (CPU.step (CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR) cpu))))) = CPU.step (CPU.Jnz CPU.REG_TEMP1 4) (CPU.step (CPU.AddConst CPU.REG_ADDR RULE_SIZE) (CPU.step (CPU.Jz CPU.REG_TEMP1 12) (CPU.step (CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q') (CPU.step (CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q) (CPU.step (CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR) cpu)))))).
  { unfold run1. rewrite Hdecode5'. reflexivity. }

  repeat split; assumption.
Qed.

(* Loop iteration lemma: checking non-matching rule preserves invariant *)
Time Lemma loop_iteration_no_match : forall tm conf cpu i,
  FindRule_Loop_Inv tm conf cpu i ->
  i < length (tm_rules tm) ->
  CPU.read_reg CPU.REG_PC cpu = 4 ->
  length cpu.(CPU.regs) = 10 ->
  decode_instr cpu = CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR ->
  decode_instr (run1 cpu) = CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q ->
  decode_instr (run_n cpu 2) =
    CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q' ->
  decode_instr (run_n cpu 3) = CPU.Jz CPU.REG_TEMP1 12 ->
  decode_instr (run_n cpu 4) = CPU.AddConst CPU.REG_ADDR RULE_SIZE ->
  decode_instr (run_n cpu 5) = CPU.Jnz CPU.REG_TEMP1 4 ->
  let '(q, tape, head) := conf in
  let sym := nth head tape (tm_blank tm) in
  let rule := nth i (tm_rules tm) (0, 0, 0, 0, 0%Z) in
  (fst (fst (fst (fst rule))), snd (fst (fst (fst rule)))) <> (q, sym) ->
  CPU.read_reg CPU.REG_TEMP1 (run_n cpu 3) <> 0 ->
  exists cpu',
    run_n cpu 6 = cpu' /\
    FindRule_Loop_Inv tm conf cpu' (S i).
Proof.
    bridge_checkpoint ("loop_iteration_no_match"%string).
Admitted.

(*
   Loop exit lemma (partial): when a matching rule is found the loop
   takes the branch into the rule payload at PC=12.  We only establish
   the first control-flow jump here; loading the rule payload and
   executing the ApplyRule block is proved separately.
 *)
Time Lemma loop_exit_match : forall tm conf cpu idx,
  FindRule_Loop_Inv tm conf cpu idx ->
  idx < length (tm_rules tm) ->
  let '(q, tape, head) := conf in
  let sym := nth head tape (tm_blank tm) in
  length cpu.(CPU.regs) = 10 ->
  decode_instr cpu = CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR ->
  decode_instr (run1 cpu) = CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q ->
  decode_instr (run_n cpu 2) =
    CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q' ->
  decode_instr (run_n cpu 3) = CPU.Jz CPU.REG_TEMP1 12 ->
  CPU.read_reg CPU.REG_TEMP1 (run_n cpu 3) = 0 ->
  exists cpu_branch,
    run_n cpu 4 = cpu_branch /\
    CPU.read_reg CPU.REG_PC cpu_branch = 12 /\
    CPU.read_reg CPU.REG_Q cpu_branch = q /\
    CPU.read_reg CPU.REG_SYM cpu_branch = sym /\
    CPU.read_reg CPU.REG_ADDR cpu_branch =
      RULES_START_ADDR + idx * RULE_SIZE.
Proof.
Admitted.

(* Main loop theorem: compose iteration lemmas *)
Time Lemma transition_FindRule_to_ApplyRule (tm : TM) (conf : TMConfig) (cpu_find : CPU.State)
  (q' write : nat) (move : Z) :
  let '(q, tape, head) := conf in
  let sym := nth head tape (tm_blank tm) in
  FindRule_Loop_Inv tm conf cpu_find 0 ->
  length cpu_find.(CPU.regs) = 10 ->
  CPU.read_reg CPU.REG_PC cpu_find = 4 ->
  decode_instr cpu_find = CPU.LoadIndirect CPU.REG_Q' CPU.REG_ADDR ->
  decode_instr (run1 cpu_find) = CPU.CopyReg CPU.REG_TEMP1 CPU.REG_Q ->
  decode_instr (run_n cpu_find 2) =
    CPU.SubReg CPU.REG_TEMP1 CPU.REG_TEMP1 CPU.REG_Q' ->
  decode_instr (run_n cpu_find 3) = CPU.Jz CPU.REG_TEMP1 12 ->
  CPU.read_reg CPU.REG_TEMP1 (run_n cpu_find 3) = 0 ->
  CPU.read_reg CPU.REG_ADDR cpu_find = RULES_START_ADDR ->
  nth 0 (tm_rules tm) (0, 0, 0, 0, 0%Z) = (q, sym, q', write, move) ->
  exists cpu_apply,
    run_n cpu_find 4 = cpu_apply /\
    CPU.read_reg CPU.REG_PC cpu_apply = 12.
Proof.
Admitted.
