(* ================================================================= *)
(* Modular Thiele Machine - Module System Variation *)
(* ================================================================= *)

(* This file is a module-based variation of the Thiele Machine.
   The MAIN WORKING IMPLEMENTATION is in ThieleMachineConcrete.v.
   
   This file has complex module system type issues between:
   - StepObs record structure
   - concrete_step predicate signature (6 arguments vs record)
   - Module signature matching requirements
   
   For the verified Thiele Machine implementation, see:
   - coq/thielemachine/coqproofs/ThieleMachineConcrete.v (WORKING)
   - coq/thielemachine/coqproofs/Subsumption.v (main theorems, PROVEN)
   - docs/FIXED_FILES_SUMMARY.md (compilation status) *)
