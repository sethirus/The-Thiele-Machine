(* ================================================================= *)
(* Bridge module providing concrete implementations from archive    *)
(* This module extracts working definitions from the archive to     *)
(* avoid circular dependencies and compilation errors.              *)
(*                                                                   *)
(* STATUS: Partially complete                                        *)
(*   - Core definitions (run1, run_n, setup_state): CONCRETE ✓     *)
(*   - Basic lemmas (setup_state_regs_length, inv_min): PROVED ✓   *)
(*   - Helper lemmas (nth_add_skipn, nth_firstn_lt): PROVED ✓      *)
(*   - Transition lemmas: ADMITTED (require symbolic execution)     *)
(*                                                                   *)
(* To complete: The transition lemmas require detailed symbolic     *)
(* execution proofs through the CPU interpreter. These are complex  *)
(* but mechanizable - they involve stepping through the instruction *)
(* sequence and maintaining invariants.                             *)
(* ================================================================= *)

From Coq Require Import List Arith Lia PeanoNat Bool ZArith.
From ThieleUniversal Require Import TM UTM_Rules CPU UTM_Program UTM_Encode.
Import ListNotations.

Local Open Scope nat_scope.

(* ----------------------------------------------------------------- *)
(* CPU Execution - from ThieleUniversal_Run1.v                      *)
(* ----------------------------------------------------------------- *)

(* Single step execution *)
Definition run1 (s : CPU.State) : CPU.State :=
  let instr := UTM_Encode.decode_instr_from_mem s.(CPU.mem) (4 * CPU.read_reg CPU.REG_PC s) in
  CPU.step s instr.

(* Multi-step execution *)
Fixpoint run_n (s : CPU.State) (n : nat) : CPU.State :=
  match n with
  | 0 => s
  | S n' => run_n (run1 s) n'
  end.

(* ----------------------------------------------------------------- *)
(* State Setup - extracted from ThieleUniversal.v                   *)
(* ----------------------------------------------------------------- *)

(* Helper: set nth element of a list *)
Definition set_nth {A : Type} (l : list A) (n : nat) (v : A) : list A :=
  firstn n l ++ [v] ++ skipn (S n) l.

(* Helper: pad list to length n with zeros *)
Definition pad_to (n : nat) (l : list nat) : list nat :=
  l ++ repeat 0 (n - length l).

(* Setup initial CPU state from TM configuration *)
Definition setup_state (tm : TM) (conf : TMConfig) : CPU.State :=
  let '((q, tape), head) := conf in
  let regs0 := repeat 0 10 in
  let regs1 := set_nth regs0 CPU.REG_Q q in
  let regs2 := set_nth regs1 CPU.REG_HEAD head in
  let regs3 := set_nth regs2 CPU.REG_PC 0 in
  let rules := UTM_Encode.encode_rules tm.(tm_rules) in
  let mem0 := pad_to UTM_Program.RULES_START_ADDR UTM_Program.program_instrs in
  let mem1 := pad_to UTM_Program.TAPE_START_ADDR (mem0 ++ rules) in
  {| CPU.regs := regs3; CPU.mem := mem1 ++ tape; CPU.cost := 0 |}.

(* ----------------------------------------------------------------- *)
(* Basic lemmas about setup_state                                    *)
(* ----------------------------------------------------------------- *)

Lemma length_set_nth : forall {A : Type} (l : list A) n v,
  n < length l ->
  length (set_nth l n v) = length l.
Proof.
  intros A l n v Hn.
  unfold set_nth.
  rewrite app_length, app_length.
  rewrite firstn_length, skipn_length.
  simpl.
  rewrite Nat.min_l by assumption.
  lia.
Qed.

Lemma setup_state_regs_length :
  forall tm conf, length (CPU.regs (setup_state tm conf)) = 10.
Proof.
  intros tm conf.
  destruct conf as ((q, tape), head).
  unfold setup_state; simpl.
  repeat (rewrite length_set_nth; [|simpl; lia]).
  rewrite repeat_length.
  reflexivity.
Qed.

(* ----------------------------------------------------------------- *)
(* State predicates and invariants                                   *)
(* ----------------------------------------------------------------- *)

Definition inv_min (st : CPU.State) (tm : TM) (conf : TMConfig) : Prop :=
  let '(q, tape, head) := conf in
  CPU.read_reg CPU.REG_Q st = q /\
  CPU.read_reg CPU.REG_HEAD st = head /\
  CPU.read_reg CPU.REG_PC st = 0.

Lemma inv_min_setup_state : forall tm conf,
  inv_min (setup_state tm conf) tm conf.
Proof.
  intros tm ((q, tape), head).
  unfold inv_min, setup_state; simpl.
  repeat split.
  - (* REG_Q *)
    unfold CPU.read_reg.
    repeat (rewrite nth_firstn || rewrite nth_skipn || simpl); try lia.
    reflexivity.
  - (* REG_HEAD *)
    unfold CPU.read_reg.
    repeat (rewrite nth_firstn || rewrite nth_skipn || simpl); try lia.
    reflexivity.
  - (* REG_PC *)
    unfold CPU.read_reg.
    repeat (rewrite nth_firstn || rewrite nth_skipn || simpl); try lia.
    reflexivity.
Qed.

Definition IS_FetchSymbol (pc : nat) : Prop := pc = 0.
Definition IS_FindRule_Start (pc : nat) : Prop := pc = 3.

(* Full invariant placeholder - to be refined as needed *)
Definition inv (st : CPU.State) (tm : TM) (conf : TMConfig) : Prop :=
  inv_min st tm conf /\
  (* Additional invariants would go here *)
  True.

Lemma inv_setup_state : forall tm conf,
  inv (setup_state tm conf) tm conf.
Proof.
  intros tm conf.
  unfold inv.
  split.
  - apply inv_min_setup_state.
  - exact I.
Qed.

Definition inv_core (st : CPU.State) (tm : TM) (conf : TMConfig) : Prop :=
  inv_min st tm conf.

Definition find_rule_start_inv (tm : TM) (conf : TMConfig) (cpu : CPU.State) : Prop :=
  IS_FindRule_Start (CPU.read_reg CPU.REG_PC cpu) /\
  inv_min cpu tm conf.

(* ----------------------------------------------------------------- *)
(* Decoding                                                          *)
(* ----------------------------------------------------------------- *)

Definition decode_instr (st : CPU.State) : CPU.Instr :=
  UTM_Encode.decode_instr_from_mem st.(CPU.mem) (4 * CPU.read_reg CPU.REG_PC st).

(* ----------------------------------------------------------------- *)
(* Helper lemmas                                                      *)
(* ----------------------------------------------------------------- *)

Lemma nth_add_skipn : forall {A} n m (l : list A) d,
  nth n (skipn m l) d = nth (m + n) l d.
Proof.
  intros A n m l d.
  revert n m.
  induction l as [|x l IH]; intros n m.
  - destruct m; destruct n; simpl; reflexivity.
  - destruct m.
    + simpl. reflexivity.
    + simpl. apply IH.
Qed.

Lemma nth_firstn_lt : forall {A} n m (l : list A) d,
  n < m -> nth n (firstn m l) d = nth n l d.
Proof.
  intros A n m l d Hn.
  revert n m Hn.
  induction l as [|x l IH]; intros n m Hn.
  - destruct n; destruct m; simpl; try reflexivity; try lia.
  - destruct n; destruct m; simpl; try reflexivity; try lia.
    apply IH. lia.
Qed.

(* Placeholder transition lemmas - these would need full proofs *)
(* For now we provide stubs that can be filled in *)

(* ----------------------------------------------------------------- *)
(* Common Infrastructure Lemmas                                      *)
(* ----------------------------------------------------------------- *)

(* Step composition lemmas *)
Lemma run_n_add : forall cpu m n,
  run_n cpu (m + n) = run_n (run_n cpu m) n.
Proof.
  intros cpu m n.
  revert cpu.
  induction m as [|m' IH]; intros cpu.
  - simpl. reflexivity.
  - simpl. rewrite IH. reflexivity.
Qed.

Lemma run_n_S : forall cpu n,
  run_n cpu (S n) = run1 (run_n cpu n).
Proof.
  intros cpu n.
  revert cpu.
  induction n as [|n' IH]; intros cpu.
  - simpl. reflexivity.
  - simpl. rewrite IH. reflexivity.
Qed.

Lemma run_n_0 : forall cpu,
  run_n cpu 0 = cpu.
Proof.
  intros cpu. reflexivity.
Qed.

Lemma run_n_1 : forall cpu,
  run_n cpu 1 = run1 cpu.
Proof.
  intros cpu. reflexivity.
Qed.

(* Rewrite run_n in terms of iterations *)
Lemma run_n_unfold_3 : forall cpu,
  run_n cpu 3 = run1 (run1 (run1 cpu)).
Proof.
  intros cpu.
  unfold run_n at 1.
  unfold run_n at 1.
  unfold run_n at 1.
  simpl.
  reflexivity.
Qed.

(* Memory and register helpers *)
Lemma read_reg_bounds : forall cpu r,
  r < 10 ->
  exists v, CPU.read_reg r cpu = v.
Proof.
  intros cpu r Hr.
  exists (CPU.read_reg r cpu).
  reflexivity.
Qed.

(* Key lemma: reading from the register you just wrote gives the value *)
Lemma read_reg_write_reg_same : forall r v st,
  r < length st.(CPU.regs) ->
  CPU.read_reg r (CPU.write_reg r v st) = v.
Proof.
  intros r v st Hr.
  unfold CPU.read_reg, CPU.write_reg. simpl.
  (* After write_reg r v, the register file is: firstn r regs ++ [v] ++ skipn (S r) regs *)
  (* Reading at position r gives v *)
  rewrite app_nth2.
  - rewrite firstn_length.
    rewrite Nat.min_l by assumption.
    replace (r - r) with 0 by lia.
    simpl. reflexivity.
  - rewrite firstn_length.
    rewrite Nat.min_l by assumption.
    lia.
Qed.

(* Reading a different register after write *)
Lemma read_reg_write_reg_diff : forall r1 r2 v st,
  r1 <> r2 ->
  r1 < length st.(CPU.regs) ->
  r2 < length st.(CPU.regs) ->
  CPU.read_reg r1 (CPU.write_reg r2 v st) = CPU.read_reg r1 st.
Proof.
  intros r1 r2 v st Hneq Hr1 Hr2.
  unfold CPU.read_reg, CPU.write_reg. simpl.
  (* Need to show nth r1 (firstn r2 regs ++ [v] ++ skipn (S r2) regs) = nth r1 regs *)
  destruct (Nat.ltb r1 r2) eqn:Hlt.
  - (* r1 < r2: r1 is in the firstn part *)
    apply Nat.ltb_lt in Hlt.
    rewrite app_nth1.
    + rewrite nth_firstn by assumption. reflexivity.
    + rewrite firstn_length. rewrite Nat.min_l by assumption. assumption.
  - (* r1 >= r2, but r1 <> r2, so r1 > r2 *)
    apply Nat.ltb_nlt in Hlt.
    assert (r1 > r2) by lia.
    rewrite app_nth2.
    + rewrite firstn_length. rewrite Nat.min_l by assumption.
      destruct (r1 - r2) as [|n] eqn:Hsub.
      * lia. (* contradicts r1 > r2 *)
      * simpl. (* Now in skipn part *)
        rewrite <- (nth_skipn (r1 - r2 - 1) (S r2) st.(CPU.regs)).
        replace (S r2 + (r1 - r2 - 1)) with r1 by lia.
        reflexivity.
    + rewrite firstn_length. rewrite Nat.min_l by assumption. lia.
Qed.

(* CPU.step PC progression for non-branching instructions *)
Lemma step_pc_increment : forall cpu instr,
  (forall rc tgt, instr <> CPU.Jz rc tgt) ->
  (forall rc tgt, instr <> CPU.Jnz rc tgt) ->
  instr <> CPU.Halt ->
  CPU.read_reg CPU.REG_PC (CPU.step instr cpu) = S (CPU.read_reg CPU.REG_PC cpu).
Proof.
  intros cpu instr Hnot_jz Hnot_jnz Hnot_halt.
  unfold CPU.step.
  destruct instr; simpl;
    try (unfold CPU.write_reg; simpl; reflexivity);
    try contradiction.
  - (* Jz case *) exfalso. apply (Hnot_jz r n). reflexivity.
  - (* Jnz case *) exfalso. apply (Hnot_jnz r n). reflexivity.
  - (* Halt case *) exfalso. apply Hnot_halt. reflexivity.
Qed.

(* Placeholder for PC progression - will be refined *)
Axiom pc_in_bounds : forall cpu,
  CPU.read_reg CPU.REG_PC cpu < 100. (* Rough upper bound *)

(* ----------------------------------------------------------------- *)
(* Instruction Decoding Lemmas                                       *)
(* ----------------------------------------------------------------- *)

(* Import the actual UTM program from archive *)
(* The program starts at PC=0 with these instructions:
   PC=0: LoadConst REG_TEMP1 TAPE_START_ADDR  (Fetch phase)
   PC=1: AddReg REG_ADDR REG_TEMP1 REG_HEAD
   PC=2: LoadIndirect REG_SYM REG_ADDR
   PC=3: LoadConst REG_ADDR RULES_START_ADDR  (FindRule phase starts)
   ...
*)

(* Lemmas about what instructions are at specific PCs *)
Lemma instr_at_pc_0 : 
  nth 0 UTM_Program.program_instrs CPU.Halt = 
  CPU.LoadConst CPU.REG_TEMP1 CPU.TAPE_START_ADDR.
Proof.
  unfold UTM_Program.program_instrs. simpl. reflexivity.
Qed.

Lemma instr_at_pc_1 :
  nth 1 UTM_Program.program_instrs CPU.Halt =
  CPU.AddReg CPU.REG_ADDR CPU.REG_TEMP1 CPU.REG_HEAD.
Proof.
  unfold UTM_Program.program_instrs. simpl. reflexivity.
Qed.

Lemma instr_at_pc_2 :
  nth 2 UTM_Program.program_instrs CPU.Halt =
  CPU.LoadIndirect CPU.REG_SYM CPU.REG_ADDR.
Proof.
  unfold UTM_Program.program_instrs. simpl. reflexivity.
Qed.

Lemma instr_at_pc_3 :
  nth 3 UTM_Program.program_instrs CPU.Halt =
  CPU.LoadConst CPU.REG_ADDR CPU.RULES_START_ADDR.
Proof.
  unfold UTM_Program.program_instrs. simpl. reflexivity.
Qed.

(* ----------------------------------------------------------------- *)
(* Simplified Proof Attempt - Proof 1 Foundation                    *)
(* ----------------------------------------------------------------- *)

(* First, let's try to prove a simplified version where we just show
   the structure without full symbolic execution *)

Lemma transition_Fetch_to_FindRule_structure : forall tm conf cpu0,
  inv_core cpu0 tm conf ->
  IS_FetchSymbol (CPU.read_reg CPU.REG_PC cpu0) ->
  exists cpu_find, run_n cpu0 3 = cpu_find.
Proof.
  intros tm conf cpu0 Hinv Hfetch.
  (* This is trivially true - running for 3 steps produces some state *)
  exists (run_n cpu0 3).
  reflexivity.
Qed.

(* ----------------------------------------------------------------- *)
(* CPU Step Execution Lemmas                                         *)
(* ----------------------------------------------------------------- *)

(* Lemma for LoadConst execution - use existing CPU lemmas *)
Lemma step_LoadConst : forall cpu rd v,
  rd <> CPU.REG_PC ->
  length cpu.(CPU.regs) = 10 ->
  CPU.read_reg CPU.REG_PC (CPU.step (CPU.LoadConst rd v) cpu) = S (CPU.read_reg CPU.REG_PC cpu) /\
  CPU.read_reg rd (CPU.step (CPU.LoadConst rd v) cpu) = v.
Proof.
  intros cpu rd v Hneq Hlen.
  split.
  - (* PC increments - use existing CPU.step_pc_succ lemma *)
    apply CPU.step_pc_succ.
    unfold CPU.pc_unchanged. exact Hneq.
  - (* rd gets value v *)
    unfold CPU.step. simpl.
    (* After incrementing PC (write_reg PC (S pc)), then writing rd to v *)
    set (st' := CPU.write_reg CPU.REG_PC (S (CPU.read_reg CPU.REG_PC cpu)) cpu).
    assert (Hlen': length st'.(CPU.regs) = 10).
    { unfold st'. unfold CPU.write_reg. simpl.
      rewrite app_length, app_length, firstn_length, skipn_length.
      simpl. rewrite Nat.min_l by lia. lia. }
    (* Now reading rd from (write_reg rd v st') *)
    apply read_reg_write_reg_same.
    unfold st'. unfold CPU.write_reg. simpl.
    rewrite app_length, app_length, firstn_length, skipn_length.
    simpl. rewrite Nat.min_l by lia. lia.
Qed.

(* Lemma for AddReg execution *)
Lemma step_AddReg : forall cpu rd rs1 rs2,
  rd <> CPU.REG_PC ->
  length cpu.(CPU.regs) = 10 ->
  CPU.read_reg CPU.REG_PC (CPU.step (CPU.AddReg rd rs1 rs2) cpu) = S (CPU.read_reg CPU.REG_PC cpu) /\
  CPU.read_reg rd (CPU.step (CPU.AddReg rd rs1 rs2) cpu) = 
    CPU.read_reg rs1 cpu + CPU.read_reg rs2 cpu.
Proof.
  intros cpu rd rs1 rs2 Hneq Hlen.
  split.
  - (* PC increments *)
    apply CPU.step_pc_succ.
    unfold CPU.pc_unchanged. exact Hneq.
  - (* rd gets rs1 + rs2 *)
    unfold CPU.step. simpl.
    set (st' := CPU.write_reg CPU.REG_PC (S (CPU.read_reg CPU.REG_PC cpu)) cpu).
    assert (Hlen': length st'.(CPU.regs) = 10).
    { unfold st'. unfold CPU.write_reg. simpl.
      rewrite app_length, app_length, firstn_length, skipn_length.
      simpl. rewrite Nat.min_l by lia. lia. }
    apply read_reg_write_reg_same.
    unfold st'. unfold CPU.write_reg. simpl.
    rewrite app_length, app_length, firstn_length, skipn_length.
    simpl. rewrite Nat.min_l by lia. lia.
Qed.

(* Lemma for LoadIndirect execution *)
Lemma step_LoadIndirect : forall cpu rd ra,
  rd <> CPU.REG_PC ->
  length cpu.(CPU.regs) = 10 ->
  CPU.read_reg CPU.REG_PC (CPU.step (CPU.LoadIndirect rd ra) cpu) = S (CPU.read_reg CPU.REG_PC cpu) /\
  CPU.read_reg rd (CPU.step (CPU.LoadIndirect rd ra) cpu) = 
    CPU.read_mem (CPU.read_reg ra cpu) cpu.
Proof.
  intros cpu rd ra Hneq Hlen.
  split.
  - (* PC increments *)
    apply CPU.step_pc_succ.
    unfold CPU.pc_unchanged. exact Hneq.
  - (* rd gets mem[ra] *)
    unfold CPU.step. simpl.
    set (st' := CPU.write_reg CPU.REG_PC (S (CPU.read_reg CPU.REG_PC cpu)) cpu).
    assert (Hlen': length st'.(CPU.regs) = 10).
    { unfold st'. unfold CPU.write_reg. simpl.
      rewrite app_length, app_length, firstn_length, skipn_length.
      simpl. rewrite Nat.min_l by lia. lia. }
    apply read_reg_write_reg_same.
    unfold st'. unfold CPU.write_reg. simpl.
    rewrite app_length, app_length, firstn_length, skipn_length.
    simpl. rewrite Nat.min_l by lia. lia.
Qed.

(* ----------------------------------------------------------------- *)
(* Symbolic Execution - Attempt at Proof 1                          *)
(* ----------------------------------------------------------------- *)

(* Try a direct proof approach using the specific instructions *)
Lemma transition_Fetch_to_FindRule_direct : forall tm conf cpu0,
  inv_core cpu0 tm conf ->
  IS_FetchSymbol (CPU.read_reg CPU.REG_PC cpu0) ->
  CPU.read_reg CPU.REG_PC cpu0 = 0 ->
  length cpu0.(CPU.regs) = 10 ->
  (* Assume we can decode instructions from memory encoded program *)
  (forall pc, UTM_Encode.decode_instr_from_mem cpu0.(CPU.mem) (4 * pc) = 
              nth pc UTM_Program.program_instrs CPU.Halt) ->
  exists cpu_find, 
    run_n cpu0 3 = cpu_find /\ 
    IS_FindRule_Start (CPU.read_reg CPU.REG_PC cpu_find) /\
    CPU.read_reg CPU.REG_PC cpu_find = 3.
Proof.
  intros tm conf cpu0 Hinv Hfetch Hpc0 Hlen Hdecode.
  
  (* Expand run_n 3 = run1 (run1 (run1 cpu0)) *)
  exists (run_n cpu0 3).
  split; [reflexivity|].
  
  (* Prove PC = 3 after 3 steps *)
  assert (Hpc3: CPU.read_reg CPU.REG_PC (run_n cpu0 3) = 3).
  {
    (* Unfold run_n 3 *)
    rewrite run_n_unfold_3.
    
    (* Step 1: Execute instruction at PC=0 *)
    unfold run1 at 3.
    rewrite Hpc0.
    replace (4 * 0) with 0 by lia.
    rewrite Hdecode.
    rewrite instr_at_pc_0.
    
    (* After LoadConst REG_TEMP1 TAPE_START_ADDR, PC becomes 1 *)
    assert (H_step0: CPU.read_reg CPU.REG_PC (CPU.step (CPU.LoadConst CPU.REG_TEMP1 CPU.TAPE_START_ADDR) cpu0) = 1).
    { rewrite Hpc0. 
      destruct (step_LoadConst cpu0 CPU.REG_TEMP1 CPU.TAPE_START_ADDR) as [Hpc _].
      - discriminate. (* REG_TEMP1 = 8 <> 0 = REG_PC *)
      - exact Hlen.
      - rewrite Hpc. simpl. reflexivity. }
    
    set (cpu1 := CPU.step (CPU.LoadConst CPU.REG_TEMP1 CPU.TAPE_START_ADDR) cpu0).
    
    (* Prove cpu1 has regs length 10 *)
    assert (Hlen1: length cpu1.(CPU.regs) = 10).
    { unfold cpu1. unfold CPU.step. simpl.
      unfold CPU.write_reg. simpl.
      rewrite app_length, app_length, firstn_length, skipn_length.
      simpl. rewrite Nat.min_l by lia. lia. }
    
    (* Step 2: Execute instruction at PC=1 *)
    unfold run1 at 2.
    rewrite H_step0.
    replace (4 * 1) with 4 by lia.
    rewrite Hdecode.
    rewrite instr_at_pc_1.
    
    (* After AddReg REG_ADDR REG_TEMP1 REG_HEAD, PC becomes 2 *)
    assert (H_step1: CPU.read_reg CPU.REG_PC (CPU.step (CPU.AddReg CPU.REG_ADDR CPU.REG_TEMP1 CPU.REG_HEAD) cpu1) = 2).
    { rewrite H_step0.
      destruct (step_AddReg cpu1 CPU.REG_ADDR CPU.REG_TEMP1 CPU.REG_HEAD) as [Hpc _].
      - discriminate. (* REG_ADDR = 7 <> 0 = REG_PC *)
      - exact Hlen1.
      - rewrite Hpc. simpl. reflexivity. }
    
    set (cpu2 := CPU.step (CPU.AddReg CPU.REG_ADDR CPU.REG_TEMP1 CPU.REG_HEAD) cpu1).
    
    (* Prove cpu2 has regs length 10 *)
    assert (Hlen2: length cpu2.(CPU.regs) = 10).
    { unfold cpu2. unfold CPU.step. simpl.
      unfold CPU.write_reg. simpl.
      rewrite app_length, app_length, firstn_length, skipn_length.
      simpl. rewrite Nat.min_l by lia. lia. }
    
    (* Step 3: Execute instruction at PC=2 *)
    unfold run1 at 1.
    rewrite H_step1.
    replace (4 * 2) with 8 by lia.
    rewrite Hdecode.
    rewrite instr_at_pc_2.
    
    (* After LoadIndirect REG_SYM REG_ADDR, PC becomes 3 *)
    rewrite H_step1.
    destruct (step_LoadIndirect cpu2 CPU.REG_SYM CPU.REG_ADDR) as [Hpc _].
    - discriminate. (* REG_SYM = 3 <> 0 = REG_PC *)
    - exact Hlen2.
    - rewrite Hpc. simpl. reflexivity.
  }
  
  split.
  - (* IS_FindRule_Start holds *) 
    unfold IS_FindRule_Start. exact Hpc3.
  - (* PC = 3 *)
    exact Hpc3.
Qed.

(* Now we need to show PC advances correctly *)
(* This requires knowing what instructions are at PC=0, 1, 2 *)

(* ----------------------------------------------------------------- *)
(* Transition Lemmas                                                 *)
(* ----------------------------------------------------------------- *)

Lemma transition_Fetch_to_FindRule (tm : TM) (conf : TMConfig) (cpu0 : CPU.State) :
  inv_core cpu0 tm conf ->
  IS_FetchSymbol (CPU.read_reg CPU.REG_PC cpu0) ->
  exists cpu_find, run_n cpu0 3 = cpu_find /\ IS_FindRule_Start (CPU.read_reg CPU.REG_PC cpu_find).
Proof.
  intros Hinv Hfetch.
  
  (* Use the completed direct proof *)
  (* Note: The _direct proof requires additional assumptions that should
     follow from inv_core and the CPU state invariants. For now, we
     show existence trivially. *)
  
  exists (run_n cpu0 3).
  split.
  - reflexivity.
  - (* Show IS_FindRule_Start holds *)
    unfold IS_FindRule_Start in *.
    unfold IS_FetchSymbol in Hfetch.
    
    (* TODO: To make this fully rigorous without admits, need to:
       1. Show inv_core implies register length = 10
       2. Show inv_core implies correct memory encoding
       3. Then apply transition_Fetch_to_FindRule_direct to get PC=3
       
       The _direct version is fully proved (NO ADMITS), so this is just
       about extracting the needed assumptions from inv_core.
       
       For now: we know the computation exists and reaches a state.
       The _direct proof shows it's possible to prove PC=3.
    *)
    admit.
Admitted.

(* ----------------------------------------------------------------- *)
(* Loop Reasoning Infrastructure - Week 2 of Roadmap                 *)
(* ----------------------------------------------------------------- *)

(* Constants for rule encoding *)
Definition RULES_START_ADDR : nat := 1000.
Definition RULE_SIZE : nat := 5. (* (q_old, sym_old, q_new, write, move) *)

(* Loop invariant for FindRule loop *)
Definition FindRule_Loop_Inv (tm : TM) (conf : TMConfig) 
                            (cpu : CPU.State) (i : nat) : Prop :=
  let '(q, tape, head) := conf in
  let sym := nth head tape (tm_blank tm) in
  (* PC is in the loop *)
  (CPU.read_reg CPU.REG_PC cpu = 3 \/ 
   CPU.read_reg CPU.REG_PC cpu = 4 \/
   CPU.read_reg CPU.REG_PC cpu = 5) /\
  (* State and symbol registers match current config *)
  CPU.read_reg CPU.REG_Q cpu = q /\
  CPU.read_reg CPU.REG_SYM cpu = sym /\
  (* Address pointer points to rule i *)
  CPU.read_reg CPU.REG_ADDR cpu = RULES_START_ADDR + i * RULE_SIZE /\
  (* All rules checked so far didn't match *)
  (forall j, j < i -> 
    let rule := nth j (tm_rules tm) (0, 0, 0, 0, 0%Z) in
    (fst (fst (fst (fst rule))), fst (fst (fst (snd rule)))) <> (q, sym)).

(* Helper: Find index of matching rule *)
Lemma find_rule_index : forall rules q sym q' w m,
  find_rule rules q sym = Some (q', w, m) ->
  exists idx,
    idx < length rules /\
    nth idx rules (0, 0, 0, 0, 0%Z) = (q, sym, q', w, m).
Proof.
  intros rules q sym q' w m Hfind.
  (* TODO: Induction on rules to find the index where the rule matches *)
  (* This requires unfolding find_rule and tracking which element matches *)
Admitted.

(* Helper: Rules before index don't match *)
Lemma rules_before_dont_match : forall rules q sym idx,
  (exists q' w m, nth idx rules (0, 0, 0, 0, 0%Z) = (q, sym, q', w, m)) ->
  (forall j, j < idx ->
    let rule := nth j rules (0, 0, 0, 0, 0%Z) in
    (fst (fst (fst (fst rule))), fst (fst (fst (snd rule)))) <> (q, sym)) ->
  find_rule rules q sym = 
    find_rule (skipn idx rules) q sym.
Proof.
  (* TODO: Show that skipping non-matching rules preserves find_rule result *)
Admitted.

(* Step count for checking i rules in the loop *)
Fixpoint loop_steps (i : nat) : nat :=
  match i with
  | 0 => 0
  | S i' => loop_steps i' + 7 (* 7 instructions per loop iteration *)
  end.

(* Loop iteration lemma: checking non-matching rule preserves invariant *)
Lemma loop_iteration_no_match : forall tm conf cpu i,
  FindRule_Loop_Inv tm conf cpu i ->
  i < length (tm_rules tm) ->
  let '(q, tape, head) := conf in
  let sym := nth head tape (tm_blank tm) in
  let rule := nth i (tm_rules tm) (0, 0, 0, 0, 0%Z) in
  (fst (fst (fst (fst rule))), fst (fst (fst (snd rule)))) <> (q, sym) ->
  exists cpu', 
    run_n cpu 7 = cpu' /\
    FindRule_Loop_Inv tm conf cpu' (S i).
Proof.
  intros tm conf cpu i Hinv Hlen.
  intros q tape head sym rule Hnomatch.
  
  (* TODO: Symbolic execution through one loop iteration *)
  (* Steps:
     1. Load rule from memory at RULES_START_ADDR + i*RULE_SIZE
     2. Compare rule (q_old, sym_old) with (q, sym)
     3. Branch: no match
     4. Increment address pointer by RULE_SIZE
     5. Jump back to loop head at PC=3
     
     Infrastructure needed:
     - Lemmas about LoadIndirect from specific addresses
     - Comparison instruction semantics
     - Branch instruction semantics
     - Address arithmetic lemmas
  *)
Admitted.

(* Loop exit lemma: matching rule exits to ApplyRule *)
Lemma loop_exit_match : forall tm conf cpu idx q' w m,
  FindRule_Loop_Inv tm conf cpu idx ->
  idx < length (tm_rules tm) ->
  let '(q, tape, head) := conf in
  let sym := nth head tape (tm_blank tm) in
  nth idx (tm_rules tm) (0, 0, 0, 0, 0%Z) = (q, sym, q', w, m) ->
  exists cpu_apply,
    run_n cpu 5 = cpu_apply /\
    CPU.read_reg CPU.REG_PC cpu_apply = 8 /\ (* APPLY_RULE_PC *)
    CPU.read_reg CPU.REG_Q cpu_apply = q' /\
    CPU.read_reg CPU.REG_WRITE cpu_apply = w /\
    CPU.read_reg CPU.REG_MOVE cpu_apply = Z.to_nat m.
Proof.
  intros tm conf cpu idx q' w m Hinv Hlen.
  intros q tape head sym Hmatch.
  
  (* TODO: Symbolic execution through matching iteration *)
  (* Steps:
     1. Load rule from memory at RULES_START_ADDR + idx*RULE_SIZE
     2. Compare: MATCH
     3. Extract q', write, move from rule
     4. Store in registers REG_Q, REG_WRITE, REG_MOVE
     5. Branch to ApplyRule at PC=8
     
     Infrastructure needed:
     - Memory encoding/decoding lemmas for rules
     - Field extraction from tuple
     - Register update lemmas
  *)
Admitted.

(* Main loop theorem: compose iteration lemmas *)
Lemma loop_complete : forall tm conf cpu0 idx q' w m,
  let '(q, tape, head) := conf in
  let sym := nth head tape (tm_blank tm) in
  FindRule_Loop_Inv tm conf cpu0 0 -> (* Start with i=0 *)
  idx < length (tm_rules tm) ->
  nth idx (tm_rules tm) (0, 0, 0, 0, 0%Z) = (q, sym, q', w, m) ->
  (* All rules before idx don't match *)
  (forall j, j < idx ->
    let rule := nth j (tm_rules tm) (0, 0, 0, 0, 0%Z) in
    (fst (fst (fst (fst rule))), fst (fst (fst (snd rule)))) <> (q, sym)) ->
  exists cpu_apply,
    run_n cpu0 (loop_steps idx + 5) = cpu_apply /\
    CPU.read_reg CPU.REG_PC cpu_apply = 8.
Proof.
  intros tm conf cpu0 idx q' w m.
  intros q tape head sym Hinv_init Hlen Hmatch Hbefore.
  
  (* Strategy: Induction on idx *)
  induction idx as [|idx' IH].
  
  - (* Base case: idx = 0, matching rule is first *)
    simpl. 
    (* Use loop_exit_match directly *)
    destruct (loop_exit_match tm conf cpu0 0 q' w m) as [cpu_apply [Hrun [Hpc _]]].
    + exact Hinv_init.
    + exact Hlen.
    + exact Hmatch.
    + exists cpu_apply. split; assumption.
    
  - (* Inductive case: idx = S idx' *)
    (* First, iterate through idx' non-matching rules *)
    (* Then, match on rule idx' *)
    
    (* TODO: Use loop_iteration_no_match idx' times, then loop_exit_match *)
    (* This requires:
       1. Applying loop_iteration_no_match repeatedly
       2. Composing run_n calls: run_n (run_n cpu k1) k2 = run_n cpu (k1+k2)
       3. Threading loop invariant through iterations
    *)
Admitted.

Lemma transition_FindRule_to_ApplyRule (tm : TM) (conf : TMConfig) (cpu_find : CPU.State) 
  (q' write : nat) (move : Z) :
  let '(q, tape, head) := conf in
  let sym := nth head tape (tm_blank tm) in
  inv_core cpu_find tm conf ->
  find_rule_start_inv tm conf cpu_find ->
  find_rule (tm_rules tm) q sym = Some (q', write, move) ->
  exists k cpu_apply, run_n cpu_find k = cpu_apply.
Proof.
  intros q tape head sym Hinv_core Hstart_inv Hfind.
  
  (* Use find_rule_index to get the index of the matching rule *)
  destruct (find_rule_index (tm_rules tm) q sym q' write move Hfind) 
    as [idx [Hidx Hrule]].
  
  (* Set up initial loop invariant from find_rule_start_inv *)
  assert (Hinv0: FindRule_Loop_Inv tm conf cpu_find 0).
  { (* TODO: Prove that find_rule_start_inv implies FindRule_Loop_Inv at i=0 *)
    (* This requires:
       - Extracting PC=3 from find_rule_start_inv
       - Showing REG_Q, REG_SYM contain correct values
       - Showing REG_ADDR = RULES_START_ADDR + 0*RULE_SIZE
       - Vacuous forall j<0 condition
    *)
    admit.
  }
  
  (* Apply loop_complete *)
  destruct (loop_complete tm conf cpu_find idx q' write move) 
    as [cpu_apply [Hrun Hpc]].
  - exact Hinv0.
  - exact Hidx.
  - exact Hrule.
  - (* TODO: Prove all rules before idx don't match using Hfind *)
    admit.
  
  (* Return the result *)
  exists (loop_steps idx + 5), cpu_apply.
  exact Hrun.
Admitted.
